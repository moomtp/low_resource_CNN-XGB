

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.types.all;

entity image_test is
    generic(TREE_RAM_BITS: positive := 13;
            NUM_CLASSES:   positive := 8;
            NUM_FEATURES:  positive := 255);
end image_test;

architecture behavior of image_test is
    
    component image
        generic(TREE_RAM_BITS: positive;
                NUM_CLASSES:   positive;
                NUM_FEATURES:  positive);
        port(-- Control signals
             Clk:   in std_logic;
             Reset: in std_logic;
             
             -- Inputs for the nodes reception (trees)
             Load_trees: in std_logic;
             Valid_node: in std_logic;
             Addr:       in std_logic_vector(TREE_RAM_BITS - 1  downto 0);
             Trees_din:  in std_logic_vector(31 downto 0);
             
             -- Inputs for the features reception (pixels)
             Load_features: in std_logic;
             Valid_feature: in std_logic;
             Features_din:  in std_logic_vector(15 downto 0);
             Last_feature:  in std_logic;
             
             -- Output signals
             --     Finish:     finish (also 'ready') signal
             --     Dout:       the selected class
             --     Greater:    the value of the selected class prediction
             --     Curr_state: the current state
             Finish:     out std_logic;
             Dout:       out std_logic_vector(log_2(NUM_CLASSES) - 1 downto 0);
             greater:    out std_logic_vector(31 downto 0);
             curr_state: out std_logic_vector(2 downto 0));
    end component;
    
    component counter is
        generic(BITS: natural);
        port(Clk:   in  std_logic;
             Reset: in  std_logic;
             Count: in  std_logic;
             Dout:  out std_logic_vector (BITS - 1 downto 0));
    end component;
    
    -- Inputs
    signal Clk:           std_logic := '0';
    signal Reset:         std_logic := '0';
    signal Load_trees:    std_logic := '0';
    signal Valid_node:    std_logic := '0';
    signal Addr:          std_logic_vector(TREE_RAM_BITS - 1 downto
                                           0) := (others => '0');
    signal Trees_din:     std_logic_vector(31 downto 0) := (others => '0');
    signal Load_features: std_logic := '0';
    signal Valid_feature: std_logic := '0';
    signal Features_din:  std_logic_vector(15 downto 0) := (others => '0');
    signal last_feature:  std_logic := '0';
    
    -- Outputs
    signal Finish:     std_logic;
    signal Dout:       std_logic_vector(log_2(NUM_CLASSES) - 1 downto 0);
    signal greater:    std_logic_vector(31 downto 0);
    signal curr_state: std_logic_vector(2 downto 0);
    
    -- Clock period definition
    constant Clk_period : time := 10 ns;
    
    -- Counter signals
    signal pc_count, hc_count: std_logic := '0';
    signal pixels, hits: std_logic_vector(15 downto 0) := (others => '0');
    
    -- Label signal
    signal class_label: std_logic_vector(log_2(NUM_CLASSES) - 1 downto 0);

begin
    
    -- Instantiate the Unit Under Test (UUT)
    uut: image
        generic map(TREE_RAM_BITS => TREE_RAM_BITS,
                    NUM_CLASSES   => NUM_CLASSES,
                    NUM_FEATURES  => NUM_FEATURES)
        port map(Clk           => Clk,
                 Reset         => Reset,
                 Load_trees    => Load_trees,
                 Valid_node    => Valid_node,
                 Addr          => Addr,
                 Trees_din     => Trees_din,
                 Load_features => Load_features,
                 Valid_feature => Valid_feature,
                 Features_din  => Features_din,
                 Last_feature  => Last_feature,
                 Finish        => Finish,
                 Dout          => Dout,
                 greater       => greater,
                 curr_state    => curr_state);
    
    -- To count the pixels
    pixel_counter: counter
        generic map(BITS => 16)
        port map(Clk   => Clk, 
                 Reset => Reset,
                 Count => pc_count,
                 Dout  => pixels);
    
    -- To count the hits
    hit_counter: counter
        generic map(BITS => 16)
        port map(Clk   => Clk, 
                 Reset => Reset,
                 Count => hc_count,
                 Dout  => hits);
    
    -- Clock process definition
    Clk_process: process
    begin
        Clk <= '0';
        wait for Clk_period/2;
        Clk <= '1';
        wait for Clk_period/2;
    end process;
    
    -- Stimulus process
    stim_proc: process
    begin
        
        Reset <= '1';
        
        -- hold reset state for 100 ns.
        wait for 100 ns;
        
        Reset <= '0';
        
        wait for Clk_period*10;
        


        
        -- LOAD TREES
        -----------------------------------------------------------------------
        
        -- Load and valid trees flags
        Load_trees <= '1';
        Valid_node <= '1';

        -- Class  0
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"12000c78";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"0b000240";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"26007e20";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"5a000410";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"1aff1b08";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"0dffcf04";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"006d01bd";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"023101bd";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"97fee404";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"fff301bd";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"033501bd";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"1b004c08";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"0700a604";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"036301bd";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"022d01bd";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"a7ff9804";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"01c001bd";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"ffbc01bd";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"f9fee010";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"0dff8608";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"1aff3604";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"ffcd01bd";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"01de01bd";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"9aff9a04";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"004601bd";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"023601bd";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"73ffd208";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"76ffeb04";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"02ff01bd";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"011101bd";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"01ff0104";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"00e601bd";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"02d101bd";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"0400461c";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"0a004c0c";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"66003608";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"03fff204";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"032901bd";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"019b01bd";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"ff7701bd";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"91fff508";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"3fffd104";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"01e601bd";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"003801bd";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"21ff8b04";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"ffa401bd";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"034901bd";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"0700020c";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"fe005908";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"0400b704";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"02b001bd";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"ffd601bd";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"ff8101bd";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"3f003208";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"5a007f04";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"fff101bd";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"017401bd";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"b4ff9b04";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"ff8101bd";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"017b01bd";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"52ff072c";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"7dff8610";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"a7ff2a04";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"02e701bd";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"eaff4704";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"014f01bd";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"05000f04";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"003701bd";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"ff6a01bd";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"07ffce0c";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"9fff6c04";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"ff7601bd";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"54ffaf04";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"ffa401bd";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"02e701bd";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"2b001b08";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"4cfeae04";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"005b01bd";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"ff5a01bd";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"49ffbe04";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"ff8201bd";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"00d801bd";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"12005d20";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"05005c10";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"4effd508";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"8a002b04";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"02ce01bd";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"002a01bd";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"d0000704";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"025501bd";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"ffeb01bd";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"0dff9b08";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"25ffbf04";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"011401bd";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"ffa901bd";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"c7fed104";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"026801bd";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"003301bd";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"07ffb40c";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"d5000304";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"032501bd";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"00ff5f04";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"003701bd";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"ffa401bd";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"e2ff6708";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"eafed204";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"012901bd";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"ff7e01bd";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"01fed504";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"ffd301bd";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"029d01bd";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"1200477c";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"0400a640";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"10fff620";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"1efeee10";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"d7005008";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"84002d04";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"01690371";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"ff730371";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"85ff9f04";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"00a10371";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"ff8c0371";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"0dff9e08";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"75009204";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"014f0371";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"002c0371";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"9aff5d04";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"01090371";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"01b10371";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"1afe3b10";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"dbffb008";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"18000604";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"ff990371";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"015d0371";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"48005204";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"ff500371";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"003c0371";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"44005308";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"a7ffb104";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"01390371";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"00770371";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"fdffaf04";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"ffb70371";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"00e50371";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"08004e1c";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"7bfebd0c";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"80ffcb04";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"ff5b0371";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"23ffb704";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"016f0371";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"ff7b0371";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"33ff3008";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"5a004504";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"ffc10371";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"01100371";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"35fedb04";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"01b00371";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"009f0371";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"b4fefb10";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"c6ff7e08";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"6effac04";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"00ab0371";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"ff830371";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"4cff3a04";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"019f0371";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"ff740371";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"98fe5908";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"afff8c04";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"ffa40371";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"02560371";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"4aff3004";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"00ac0371";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"ff570371";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"d700372c";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"52ff2910";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"29ff0008";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"24ff8004";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"01530371";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"00320371";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"deff0a04";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"003d0371";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"ff630371";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"f0ff0a0c";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"bfff9f08";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"b4fe6404";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"003b0371";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"ff6f0371";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"01a70371";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"1b002708";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"f8008404";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"023b0371";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"002e0371";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"35fee904";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"ff8b0371";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"01430371";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"7efecf18";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"52ffc210";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"5a00f308";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"6eff7504";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"00180371";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"ff550371";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"3fffda04";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"01490371";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"ff770371";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"34001e04";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"01a00371";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"ffa10371";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"37ffd410";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"1bff9608";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"b3ff3f04";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"ffc20371";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"01df0371";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"8b007804";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"ff650371";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"01350371";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"16ff1e08";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"16fe7d04";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"009e0371";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"02450371";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"ffa80371";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"53001f7c";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"04009540";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"7d002720";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"d7007410";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"09000008";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"11001704";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"012304e5";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"ffa504e5";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"2bfef904";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"ffb604e5";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"00d504e5";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"e9fe4e08";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"91ffdb04";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"ffb304e5";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"00a204e5";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"21ffdf04";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"009a04e5";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"011c04e5";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"04000410";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"26004508";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"0a00f304";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"014904e5";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"ff8204e5";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"91ff7e04";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"ffa104e5";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"00c304e5";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"5a007108";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"e1ff5904";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"00be04e5";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"ffad04e5";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"1b000204";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"00c204e5";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"ffc904e5";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"07008b20";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"3f004310";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"de002408";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"9cff7b04";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"00e504e5";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"001504e5";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"09008104";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"015904e5";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"ff8704e5";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"fdffb108";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"9fff1a04";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"ff5204e5";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"001f04e5";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"d1ff3204";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"010e04e5";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"ffd804e5";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"4fffb310";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"6cff9408";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"00ff1c04";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"008404e5";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"ff6f04e5";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"7efeb504";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"fffd04e5";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"013204e5";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"61ff9504";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"ff5704e5";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"1afedc04";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"ff7104e5";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"011104e5";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"0dff3818";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"57ffe010";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"12ff5a04";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"005f04e5";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"c3009f08";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"1aff5304";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"ff5504e5";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"000504e5";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"003704e5";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"0a007804";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"015b04e5";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"ffaa04e5";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"5a00e21c";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"5fffaa10";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"d5ff8408";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"67ff3904";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"016d04e5";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"001c04e5";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"52ff8804";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"ff7704e5";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"006804e5";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"8fff2b08";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"97fe9204";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"002b04e5";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"01a804e5";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"ff7904e5";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"08005508";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"78ffe704";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"019204e5";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"fffe04e5";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"ff6f04e5";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"fe003070";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"75009e40";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"2bff4320";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"76ffa410";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"b6ff7408";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"5100a404";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"00e80649";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"ff960649";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"22ffe804";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"ff690649";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"00650649";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"10ffd508";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"25004404";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"00780649";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"ffae0649";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"75ff6a04";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"00bd0649";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"ff940649";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"93ff7f10";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"fafe9708";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"adffa804";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"ff610649";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"01110649";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"4e004804";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"00d40649";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"ffd10649";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"62ff5d08";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"7dffef04";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"00880649";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"00070649";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"3eff8904";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"00e30649";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"00660649";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"0dffb018";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"1dfef70c";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"93ffca08";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"40ffe104";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"ffc00649";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"01340649";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"ff630649";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"e2ffef08";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"d2fe5c04";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"00510649";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"ff5c0649";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"01240649";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"b2ffd20c";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"bfffbd04";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"ff480649";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"04fffe04";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"00ca0649";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"fff80649";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"8a002408";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"66004d04";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"01020649";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"ffc10649";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"ff660649";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"26003924";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"24ffa710";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"d5fff50c";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"9bff2b04";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"ff660649";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"7aff8104";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"014a0649";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"fff50649";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"ff560649";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"99fe6804";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"ff6a0649";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"40ffbd08";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"24ffec04";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"00270649";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"ff750649";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"ebfe9304";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"ff9a0649";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"01390649";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"0affb510";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"7dffb408";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"36ffa404";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"015c0649";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"ffa20649";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"27ff4d04";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"00390649";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"ff620649";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"0cfd6b04";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"00b10649";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"38007f08";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"de00b304";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"ff670649";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"003f0649";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"00b30649";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"52ff0364";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"0dff6d38";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"76ffec20";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"08006110";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"65ff3f08";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"feffc904";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"007007e5";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"ff6807e5";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"27ffba04";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"011107e5";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"002807e5";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"e1ff0a08";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"03ff8804";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"011607e5";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"001207e5";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"c6ff1d04";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"ff5f07e5";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"ffe907e5";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"7eff5410";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"f6ffa708";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"75ff0a04";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"00be07e5";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"ff6807e5";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"71ff4404";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"ff9107e5";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"011a07e5";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"8efffa04";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"ff8b07e5";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"012807e5";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"33fef914";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"f9ffe310";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"e4ff1b08";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"7ffdee04";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"00fb07e5";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"ff5807e5";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"44000804";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"011407e5";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"ff9707e5";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"00db07e5";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"4effed10";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"31005208";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"c2fff904";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"00b807e5";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"ff9507e5";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"8b000804";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"ff7d07e5";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"007607e5";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"07009804";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"ff4e07e5";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"002b07e5";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"4cffb040";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"3f004a20";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"43ff4110";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"63ffce08";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"baff8c04";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"003507e5";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"009b07e5";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"f5002f04";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"ffba07e5";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"009707e5";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"11001d08";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"e9fe3a04";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"004c07e5";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"00b507e5";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"01fef304";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"ff5207e5";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"00ae07e5";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"08008410";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"55008008";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"6a000c04";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"005307e5";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"ff8007e5";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"0dfeff04";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"ff6307e5";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"00e707e5";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"20ff6e08";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"7bfef404";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"ff7c07e5";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"009d07e5";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"27ff9a04";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"001b07e5";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"ff4207e5";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"07ffc20c";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"7efe2504";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"ff8a07e5";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"25ffc304";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"000307e5";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"011d07e5";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"cdffea10";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"daff4608";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"46feb204";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"ff7307e5";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"00d107e5";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"65001a04";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"ff6707e5";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"00b307e5";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"10ffbe08";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"89002004";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"00cd07e5";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"ff8707e5";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"f5005404";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"ff8107e5";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"00c807e5";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"12005d70";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"4efff240";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"3100b620";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"63ffd610";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"40001108";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"52fe8304";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"ff9c0939";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"00930939";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"65ff3604";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"00220939";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"00740939";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"6affd808";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"deffa204";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"ffc20939";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"00730939";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"31fef604";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"00b60939";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"ffcb0939";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"37ff9410";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"4bfe3008";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"8b003d04";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"ff990939";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"00f30939";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"54001e04";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"00080939";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"ff450939";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"9affab08";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"46ff9704";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"ff4c0939";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"00740939";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"cc007304";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"00da0939";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"ff6a0939";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"bfff741c";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"59003f10";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"9dff7a08";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"1e005804";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"ffa40939";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"01050939";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"c7ffc104";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"ff460939";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"00740939";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"d6008d08";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"d3fe9704";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"fff40939";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"010e0939";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"ff5e0939";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"44007510";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"9bff6408";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"a7ffed04";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"003e0939";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"ff630939";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"d4ff1d04";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"ffb30939";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"00df0939";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"ff420939";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"37ffdb24";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"0dffcc18";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"63ff0508";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"fdfef104";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"00d70939";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"ff960939";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"5a00f308";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"0aff7d04";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"00680939";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"ff620939";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"33ff1804";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"ff870939";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"009d0939";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"a5feb404";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"01020939";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"67ffe904";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"ff690939";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"00ba0939";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"7efea908";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"17004504";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"ff620939";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"00a30939";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"5effa104";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"ff990939";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"b9fe4e04";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"00000939";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"77ff8004";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"01140939";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"004a0939";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"fe002a80";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"4fff6140";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"21ffe320";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"e3fe5010";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"28ff4308";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"eaff7f04";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"ff520acd";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"fffe0acd";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"3eff9f04";
		wait for Clk_period;
		Addr <=  "0001001010111";
		Trees_din <= x"00650acd";
		wait for Clk_period;
		Addr <=  "0001001011000";
		Trees_din <= x"ff910acd";
		wait for Clk_period;
		Addr <=  "0001001011001";
		Trees_din <= x"d5009d08";
		wait for Clk_period;
		Addr <=  "0001001011010";
		Trees_din <= x"7dff7504";
		wait for Clk_period;
		Addr <=  "0001001011011";
		Trees_din <= x"008b0acd";
		wait for Clk_period;
		Addr <=  "0001001011100";
		Trees_din <= x"00470acd";
		wait for Clk_period;
		Addr <=  "0001001011101";
		Trees_din <= x"78fee004";
		wait for Clk_period;
		Addr <=  "0001001011110";
		Trees_din <= x"008f0acd";
		wait for Clk_period;
		Addr <=  "0001001011111";
		Trees_din <= x"ff400acd";
		wait for Clk_period;
		Addr <=  "0001001100000";
		Trees_din <= x"60fff110";
		wait for Clk_period;
		Addr <=  "0001001100001";
		Trees_din <= x"fafe9708";
		wait for Clk_period;
		Addr <=  "0001001100010";
		Trees_din <= x"a3ff1704";
		wait for Clk_period;
		Addr <=  "0001001100011";
		Trees_din <= x"00430acd";
		wait for Clk_period;
		Addr <=  "0001001100100";
		Trees_din <= x"ff120acd";
		wait for Clk_period;
		Addr <=  "0001001100101";
		Trees_din <= x"0cff5604";
		wait for Clk_period;
		Addr <=  "0001001100110";
		Trees_din <= x"00a60acd";
		wait for Clk_period;
		Addr <=  "0001001100111";
		Trees_din <= x"fff10acd";
		wait for Clk_period;
		Addr <=  "0001001101000";
		Trees_din <= x"b3ff3308";
		wait for Clk_period;
		Addr <=  "0001001101001";
		Trees_din <= x"aa000104";
		wait for Clk_period;
		Addr <=  "0001001101010";
		Trees_din <= x"00a50acd";
		wait for Clk_period;
		Addr <=  "0001001101011";
		Trees_din <= x"ff4a0acd";
		wait for Clk_period;
		Addr <=  "0001001101100";
		Trees_din <= x"c9ff8a04";
		wait for Clk_period;
		Addr <=  "0001001101101";
		Trees_din <= x"00570acd";
		wait for Clk_period;
		Addr <=  "0001001101110";
		Trees_din <= x"ff240acd";
		wait for Clk_period;
		Addr <=  "0001001101111";
		Trees_din <= x"87ff7720";
		wait for Clk_period;
		Addr <=  "0001001110000";
		Trees_din <= x"75008b10";
		wait for Clk_period;
		Addr <=  "0001001110001";
		Trees_din <= x"20ff6c08";
		wait for Clk_period;
		Addr <=  "0001001110010";
		Trees_din <= x"da004104";
		wait for Clk_period;
		Addr <=  "0001001110011";
		Trees_din <= x"006a0acd";
		wait for Clk_period;
		Addr <=  "0001001110100";
		Trees_din <= x"ffbe0acd";
		wait for Clk_period;
		Addr <=  "0001001110101";
		Trees_din <= x"b0ff2304";
		wait for Clk_period;
		Addr <=  "0001001110110";
		Trees_din <= x"ff9d0acd";
		wait for Clk_period;
		Addr <=  "0001001110111";
		Trees_din <= x"00140acd";
		wait for Clk_period;
		Addr <=  "0001001111000";
		Trees_din <= x"d7ffff08";
		wait for Clk_period;
		Addr <=  "0001001111001";
		Trees_din <= x"6d005c04";
		wait for Clk_period;
		Addr <=  "0001001111010";
		Trees_din <= x"00c10acd";
		wait for Clk_period;
		Addr <=  "0001001111011";
		Trees_din <= x"ff6e0acd";
		wait for Clk_period;
		Addr <=  "0001001111100";
		Trees_din <= x"0bffbd04";
		wait for Clk_period;
		Addr <=  "0001001111101";
		Trees_din <= x"fff90acd";
		wait for Clk_period;
		Addr <=  "0001001111110";
		Trees_din <= x"ff6f0acd";
		wait for Clk_period;
		Addr <=  "0001001111111";
		Trees_din <= x"06ff8f10";
		wait for Clk_period;
		Addr <=  "0001010000000";
		Trees_din <= x"20ff7108";
		wait for Clk_period;
		Addr <=  "0001010000001";
		Trees_din <= x"60ffe304";
		wait for Clk_period;
		Addr <=  "0001010000010";
		Trees_din <= x"008e0acd";
		wait for Clk_period;
		Addr <=  "0001010000011";
		Trees_din <= x"ff3a0acd";
		wait for Clk_period;
		Addr <=  "0001010000100";
		Trees_din <= x"b4ff8e04";
		wait for Clk_period;
		Addr <=  "0001010000101";
		Trees_din <= x"ffcc0acd";
		wait for Clk_period;
		Addr <=  "0001010000110";
		Trees_din <= x"006a0acd";
		wait for Clk_period;
		Addr <=  "0001010000111";
		Trees_din <= x"3eff8408";
		wait for Clk_period;
		Addr <=  "0001010001000";
		Trees_din <= x"5400ce04";
		wait for Clk_period;
		Addr <=  "0001010001001";
		Trees_din <= x"00b60acd";
		wait for Clk_period;
		Addr <=  "0001010001010";
		Trees_din <= x"ffae0acd";
		wait for Clk_period;
		Addr <=  "0001010001011";
		Trees_din <= x"f1ff6d04";
		wait for Clk_period;
		Addr <=  "0001010001100";
		Trees_din <= x"ffba0acd";
		wait for Clk_period;
		Addr <=  "0001010001101";
		Trees_din <= x"00680acd";
		wait for Clk_period;
		Addr <=  "0001010001110";
		Trees_din <= x"d8004c2c";
		wait for Clk_period;
		Addr <=  "0001010001111";
		Trees_din <= x"0700601c";
		wait for Clk_period;
		Addr <=  "0001010010000";
		Trees_din <= x"b3fed40c";
		wait for Clk_period;
		Addr <=  "0001010010001";
		Trees_din <= x"29ff5a04";
		wait for Clk_period;
		Addr <=  "0001010010010";
		Trees_din <= x"ff4f0acd";
		wait for Clk_period;
		Addr <=  "0001010010011";
		Trees_din <= x"52ff3204";
		wait for Clk_period;
		Addr <=  "0001010010100";
		Trees_din <= x"ff780acd";
		wait for Clk_period;
		Addr <=  "0001010010101";
		Trees_din <= x"00c30acd";
		wait for Clk_period;
		Addr <=  "0001010010110";
		Trees_din <= x"5a003e08";
		wait for Clk_period;
		Addr <=  "0001010010111";
		Trees_din <= x"d7006404";
		wait for Clk_period;
		Addr <=  "0001010011000";
		Trees_din <= x"ff730acd";
		wait for Clk_period;
		Addr <=  "0001010011001";
		Trees_din <= x"00660acd";
		wait for Clk_period;
		Addr <=  "0001010011010";
		Trees_din <= x"a4fff304";
		wait for Clk_period;
		Addr <=  "0001010011011";
		Trees_din <= x"00d70acd";
		wait for Clk_period;
		Addr <=  "0001010011100";
		Trees_din <= x"ff7a0acd";
		wait for Clk_period;
		Addr <=  "0001010011101";
		Trees_din <= x"69ff7e04";
		wait for Clk_period;
		Addr <=  "0001010011110";
		Trees_din <= x"ff580acd";
		wait for Clk_period;
		Addr <=  "0001010011111";
		Trees_din <= x"2bff7004";
		wait for Clk_period;
		Addr <=  "0001010100000";
		Trees_din <= x"ff780acd";
		wait for Clk_period;
		Addr <=  "0001010100001";
		Trees_din <= x"64ff2a04";
		wait for Clk_period;
		Addr <=  "0001010100010";
		Trees_din <= x"00020acd";
		wait for Clk_period;
		Addr <=  "0001010100011";
		Trees_din <= x"010d0acd";
		wait for Clk_period;
		Addr <=  "0001010100100";
		Trees_din <= x"5a010714";
		wait for Clk_period;
		Addr <=  "0001010100101";
		Trees_din <= x"e000030c";
		wait for Clk_period;
		Addr <=  "0001010100110";
		Trees_din <= x"92005708";
		wait for Clk_period;
		Addr <=  "0001010100111";
		Trees_din <= x"ea007504";
		wait for Clk_period;
		Addr <=  "0001010101000";
		Trees_din <= x"ff4d0acd";
		wait for Clk_period;
		Addr <=  "0001010101001";
		Trees_din <= x"002f0acd";
		wait for Clk_period;
		Addr <=  "0001010101010";
		Trees_din <= x"003c0acd";
		wait for Clk_period;
		Addr <=  "0001010101011";
		Trees_din <= x"0affb004";
		wait for Clk_period;
		Addr <=  "0001010101100";
		Trees_din <= x"00ca0acd";
		wait for Clk_period;
		Addr <=  "0001010101101";
		Trees_din <= x"ff8f0acd";
		wait for Clk_period;
		Addr <=  "0001010101110";
		Trees_din <= x"59ff9008";
		wait for Clk_period;
		Addr <=  "0001010101111";
		Trees_din <= x"08000c04";
		wait for Clk_period;
		Addr <=  "0001010110000";
		Trees_din <= x"008c0acd";
		wait for Clk_period;
		Addr <=  "0001010110001";
		Trees_din <= x"ff640acd";
		wait for Clk_period;
		Addr <=  "0001010110010";
		Trees_din <= x"00c70acd";
		wait for Clk_period;
		Addr <=  "0001010110011";
		Trees_din <= x"0dff9e78";
		wait for Clk_period;
		Addr <=  "0001010110100";
		Trees_din <= x"52fece38";
		wait for Clk_period;
		Addr <=  "0001010110101";
		Trees_din <= x"c8ffd320";
		wait for Clk_period;
		Addr <=  "0001010110110";
		Trees_din <= x"cbffbf10";
		wait for Clk_period;
		Addr <=  "0001010110111";
		Trees_din <= x"4cff7e08";
		wait for Clk_period;
		Addr <=  "0001010111000";
		Trees_din <= x"40006b04";
		wait for Clk_period;
		Addr <=  "0001010111001";
		Trees_din <= x"00e40c89";
		wait for Clk_period;
		Addr <=  "0001010111010";
		Trees_din <= x"ff880c89";
		wait for Clk_period;
		Addr <=  "0001010111011";
		Trees_din <= x"aaff4f04";
		wait for Clk_period;
		Addr <=  "0001010111100";
		Trees_din <= x"001f0c89";
		wait for Clk_period;
		Addr <=  "0001010111101";
		Trees_din <= x"ff710c89";
		wait for Clk_period;
		Addr <=  "0001010111110";
		Trees_din <= x"26002a08";
		wait for Clk_period;
		Addr <=  "0001010111111";
		Trees_din <= x"45fe6504";
		wait for Clk_period;
		Addr <=  "0001011000000";
		Trees_din <= x"ffa50c89";
		wait for Clk_period;
		Addr <=  "0001011000001";
		Trees_din <= x"00a20c89";
		wait for Clk_period;
		Addr <=  "0001011000010";
		Trees_din <= x"89010604";
		wait for Clk_period;
		Addr <=  "0001011000011";
		Trees_din <= x"ff570c89";
		wait for Clk_period;
		Addr <=  "0001011000100";
		Trees_din <= x"001e0c89";
		wait for Clk_period;
		Addr <=  "0001011000101";
		Trees_din <= x"44ff4a08";
		wait for Clk_period;
		Addr <=  "0001011000110";
		Trees_din <= x"65ff8404";
		wait for Clk_period;
		Addr <=  "0001011000111";
		Trees_din <= x"ff9c0c89";
		wait for Clk_period;
		Addr <=  "0001011001000";
		Trees_din <= x"00f10c89";
		wait for Clk_period;
		Addr <=  "0001011001001";
		Trees_din <= x"7eff6108";
		wait for Clk_period;
		Addr <=  "0001011001010";
		Trees_din <= x"4cfe8b04";
		wait for Clk_period;
		Addr <=  "0001011001011";
		Trees_din <= x"00380c89";
		wait for Clk_period;
		Addr <=  "0001011001100";
		Trees_din <= x"ff6a0c89";
		wait for Clk_period;
		Addr <=  "0001011001101";
		Trees_din <= x"95ff6304";
		wait for Clk_period;
		Addr <=  "0001011001110";
		Trees_din <= x"ff990c89";
		wait for Clk_period;
		Addr <=  "0001011001111";
		Trees_din <= x"00aa0c89";
		wait for Clk_period;
		Addr <=  "0001011010000";
		Trees_din <= x"c2ff8b20";
		wait for Clk_period;
		Addr <=  "0001011010001";
		Trees_din <= x"3f005010";
		wait for Clk_period;
		Addr <=  "0001011010010";
		Trees_din <= x"1b006a08";
		wait for Clk_period;
		Addr <=  "0001011010011";
		Trees_din <= x"ddfef604";
		wait for Clk_period;
		Addr <=  "0001011010100";
		Trees_din <= x"00210c89";
		wait for Clk_period;
		Addr <=  "0001011010101";
		Trees_din <= x"00640c89";
		wait for Clk_period;
		Addr <=  "0001011010110";
		Trees_din <= x"1cff2e04";
		wait for Clk_period;
		Addr <=  "0001011010111";
		Trees_din <= x"00720c89";
		wait for Clk_period;
		Addr <=  "0001011011000";
		Trees_din <= x"ff5c0c89";
		wait for Clk_period;
		Addr <=  "0001011011001";
		Trees_din <= x"3aff2508";
		wait for Clk_period;
		Addr <=  "0001011011010";
		Trees_din <= x"bd005f04";
		wait for Clk_period;
		Addr <=  "0001011011011";
		Trees_din <= x"ff650c89";
		wait for Clk_period;
		Addr <=  "0001011011100";
		Trees_din <= x"00440c89";
		wait for Clk_period;
		Addr <=  "0001011011101";
		Trees_din <= x"55ffb604";
		wait for Clk_period;
		Addr <=  "0001011011110";
		Trees_din <= x"ff990c89";
		wait for Clk_period;
		Addr <=  "0001011011111";
		Trees_din <= x"003d0c89";
		wait for Clk_period;
		Addr <=  "0001011100000";
		Trees_din <= x"72006a10";
		wait for Clk_period;
		Addr <=  "0001011100001";
		Trees_din <= x"da001008";
		wait for Clk_period;
		Addr <=  "0001011100010";
		Trees_din <= x"3d001304";
		wait for Clk_period;
		Addr <=  "0001011100011";
		Trees_din <= x"ffef0c89";
		wait for Clk_period;
		Addr <=  "0001011100100";
		Trees_din <= x"00820c89";
		wait for Clk_period;
		Addr <=  "0001011100101";
		Trees_din <= x"f9fff704";
		wait for Clk_period;
		Addr <=  "0001011100110";
		Trees_din <= x"ff9e0c89";
		wait for Clk_period;
		Addr <=  "0001011100111";
		Trees_din <= x"00c80c89";
		wait for Clk_period;
		Addr <=  "0001011101000";
		Trees_din <= x"c2ff9208";
		wait for Clk_period;
		Addr <=  "0001011101001";
		Trees_din <= x"b0ff5d04";
		wait for Clk_period;
		Addr <=  "0001011101010";
		Trees_din <= x"ffdb0c89";
		wait for Clk_period;
		Addr <=  "0001011101011";
		Trees_din <= x"00c40c89";
		wait for Clk_period;
		Addr <=  "0001011101100";
		Trees_din <= x"aeffab04";
		wait for Clk_period;
		Addr <=  "0001011101101";
		Trees_din <= x"ff3d0c89";
		wait for Clk_period;
		Addr <=  "0001011101110";
		Trees_din <= x"00400c89";
		wait for Clk_period;
		Addr <=  "0001011101111";
		Trees_din <= x"4cff062c";
		wait for Clk_period;
		Addr <=  "0001011110000";
		Trees_din <= x"fafe970c";
		wait for Clk_period;
		Addr <=  "0001011110001";
		Trees_din <= x"6cff2c04";
		wait for Clk_period;
		Addr <=  "0001011110010";
		Trees_din <= x"00760c89";
		wait for Clk_period;
		Addr <=  "0001011110011";
		Trees_din <= x"32fe7b04";
		wait for Clk_period;
		Addr <=  "0001011110100";
		Trees_din <= x"ffe60c89";
		wait for Clk_period;
		Addr <=  "0001011110101";
		Trees_din <= x"ff190c89";
		wait for Clk_period;
		Addr <=  "0001011110110";
		Trees_din <= x"0800c810";
		wait for Clk_period;
		Addr <=  "0001011110111";
		Trees_din <= x"6a001c08";
		wait for Clk_period;
		Addr <=  "0001011111000";
		Trees_din <= x"90ff7404";
		wait for Clk_period;
		Addr <=  "0001011111001";
		Trees_din <= x"009b0c89";
		wait for Clk_period;
		Addr <=  "0001011111010";
		Trees_din <= x"00530c89";
		wait for Clk_period;
		Addr <=  "0001011111011";
		Trees_din <= x"ebff1804";
		wait for Clk_period;
		Addr <=  "0001011111100";
		Trees_din <= x"ffaa0c89";
		wait for Clk_period;
		Addr <=  "0001011111101";
		Trees_din <= x"00cb0c89";
		wait for Clk_period;
		Addr <=  "0001011111110";
		Trees_din <= x"76ff5b08";
		wait for Clk_period;
		Addr <=  "0001011111111";
		Trees_din <= x"a9ff0904";
		wait for Clk_period;
		Addr <=  "0001100000000";
		Trees_din <= x"00650c89";
		wait for Clk_period;
		Addr <=  "0001100000001";
		Trees_din <= x"ff310c89";
		wait for Clk_period;
		Addr <=  "0001100000010";
		Trees_din <= x"9bff3704";
		wait for Clk_period;
		Addr <=  "0001100000011";
		Trees_din <= x"ffe00c89";
		wait for Clk_period;
		Addr <=  "0001100000100";
		Trees_din <= x"00940c89";
		wait for Clk_period;
		Addr <=  "0001100000101";
		Trees_din <= x"7d002620";
		wait for Clk_period;
		Addr <=  "0001100000110";
		Trees_din <= x"10fff310";
		wait for Clk_period;
		Addr <=  "0001100000111";
		Trees_din <= x"9bfeda08";
		wait for Clk_period;
		Addr <=  "0001100001000";
		Trees_din <= x"78ff7404";
		wait for Clk_period;
		Addr <=  "0001100001001";
		Trees_din <= x"ff7a0c89";
		wait for Clk_period;
		Addr <=  "0001100001010";
		Trees_din <= x"00510c89";
		wait for Clk_period;
		Addr <=  "0001100001011";
		Trees_din <= x"95feb704";
		wait for Clk_period;
		Addr <=  "0001100001100";
		Trees_din <= x"000f0c89";
		wait for Clk_period;
		Addr <=  "0001100001101";
		Trees_din <= x"00800c89";
		wait for Clk_period;
		Addr <=  "0001100001110";
		Trees_din <= x"11fefa08";
		wait for Clk_period;
		Addr <=  "0001100001111";
		Trees_din <= x"81ffbf04";
		wait for Clk_period;
		Addr <=  "0001100010000";
		Trees_din <= x"00e70c89";
		wait for Clk_period;
		Addr <=  "0001100010001";
		Trees_din <= x"ff810c89";
		wait for Clk_period;
		Addr <=  "0001100010010";
		Trees_din <= x"77fee104";
		wait for Clk_period;
		Addr <=  "0001100010011";
		Trees_din <= x"ff730c89";
		wait for Clk_period;
		Addr <=  "0001100010100";
		Trees_din <= x"000d0c89";
		wait for Clk_period;
		Addr <=  "0001100010101";
		Trees_din <= x"ddfed40c";
		wait for Clk_period;
		Addr <=  "0001100010110";
		Trees_din <= x"8dfd5b04";
		wait for Clk_period;
		Addr <=  "0001100010111";
		Trees_din <= x"004e0c89";
		wait for Clk_period;
		Addr <=  "0001100011000";
		Trees_din <= x"8dfef004";
		wait for Clk_period;
		Addr <=  "0001100011001";
		Trees_din <= x"ff240c89";
		wait for Clk_period;
		Addr <=  "0001100011010";
		Trees_din <= x"00020c89";
		wait for Clk_period;
		Addr <=  "0001100011011";
		Trees_din <= x"12ffe208";
		wait for Clk_period;
		Addr <=  "0001100011100";
		Trees_din <= x"cf008a04";
		wait for Clk_period;
		Addr <=  "0001100011101";
		Trees_din <= x"009a0c89";
		wait for Clk_period;
		Addr <=  "0001100011110";
		Trees_din <= x"ff510c89";
		wait for Clk_period;
		Addr <=  "0001100011111";
		Trees_din <= x"87ff7004";
		wait for Clk_period;
		Addr <=  "0001100100000";
		Trees_din <= x"ff490c89";
		wait for Clk_period;
		Addr <=  "0001100100001";
		Trees_din <= x"00260c89";
		wait for Clk_period;
		Addr <=  "0001100100010";
		Trees_din <= x"93ff7e78";
		wait for Clk_period;
		Addr <=  "0001100100011";
		Trees_din <= x"1aff3840";
		wait for Clk_period;
		Addr <=  "0001100100100";
		Trees_din <= x"5d001a20";
		wait for Clk_period;
		Addr <=  "0001100100101";
		Trees_din <= x"dc003e10";
		wait for Clk_period;
		Addr <=  "0001100100110";
		Trees_din <= x"c9005c08";
		wait for Clk_period;
		Addr <=  "0001100100111";
		Trees_din <= x"80ffa304";
		wait for Clk_period;
		Addr <=  "0001100101000";
		Trees_din <= x"004a0e65";
		wait for Clk_period;
		Addr <=  "0001100101001";
		Trees_din <= x"000d0e65";
		wait for Clk_period;
		Addr <=  "0001100101010";
		Trees_din <= x"97ff9e04";
		wait for Clk_period;
		Addr <=  "0001100101011";
		Trees_din <= x"ff490e65";
		wait for Clk_period;
		Addr <=  "0001100101100";
		Trees_din <= x"00900e65";
		wait for Clk_period;
		Addr <=  "0001100101101";
		Trees_din <= x"08004608";
		wait for Clk_period;
		Addr <=  "0001100101110";
		Trees_din <= x"84fffe04";
		wait for Clk_period;
		Addr <=  "0001100101111";
		Trees_din <= x"005b0e65";
		wait for Clk_period;
		Addr <=  "0001100110000";
		Trees_din <= x"ff770e65";
		wait for Clk_period;
		Addr <=  "0001100110001";
		Trees_din <= x"58ff3a04";
		wait for Clk_period;
		Addr <=  "0001100110010";
		Trees_din <= x"ff4b0e65";
		wait for Clk_period;
		Addr <=  "0001100110011";
		Trees_din <= x"00020e65";
		wait for Clk_period;
		Addr <=  "0001100110100";
		Trees_din <= x"f8fff310";
		wait for Clk_period;
		Addr <=  "0001100110101";
		Trees_din <= x"4bfe8a08";
		wait for Clk_period;
		Addr <=  "0001100110110";
		Trees_din <= x"37ff5204";
		wait for Clk_period;
		Addr <=  "0001100110111";
		Trees_din <= x"ffff0e65";
		wait for Clk_period;
		Addr <=  "0001100111000";
		Trees_din <= x"00c30e65";
		wait for Clk_period;
		Addr <=  "0001100111001";
		Trees_din <= x"a7ff0604";
		wait for Clk_period;
		Addr <=  "0001100111010";
		Trees_din <= x"008f0e65";
		wait for Clk_period;
		Addr <=  "0001100111011";
		Trees_din <= x"ff610e65";
		wait for Clk_period;
		Addr <=  "0001100111100";
		Trees_din <= x"0400bf08";
		wait for Clk_period;
		Addr <=  "0001100111101";
		Trees_din <= x"d2ff9304";
		wait for Clk_period;
		Addr <=  "0001100111110";
		Trees_din <= x"00a90e65";
		wait for Clk_period;
		Addr <=  "0001100111111";
		Trees_din <= x"ff6f0e65";
		wait for Clk_period;
		Addr <=  "0001101000000";
		Trees_din <= x"cd000604";
		wait for Clk_period;
		Addr <=  "0001101000001";
		Trees_din <= x"ff5e0e65";
		wait for Clk_period;
		Addr <=  "0001101000010";
		Trees_din <= x"00770e65";
		wait for Clk_period;
		Addr <=  "0001101000011";
		Trees_din <= x"75005220";
		wait for Clk_period;
		Addr <=  "0001101000100";
		Trees_din <= x"c0ff2d10";
		wait for Clk_period;
		Addr <=  "0001101000101";
		Trees_din <= x"64ff0708";
		wait for Clk_period;
		Addr <=  "0001101000110";
		Trees_din <= x"f0fec704";
		wait for Clk_period;
		Addr <=  "0001101000111";
		Trees_din <= x"ffe10e65";
		wait for Clk_period;
		Addr <=  "0001101001000";
		Trees_din <= x"00ca0e65";
		wait for Clk_period;
		Addr <=  "0001101001001";
		Trees_din <= x"68feac04";
		wait for Clk_period;
		Addr <=  "0001101001010";
		Trees_din <= x"ff910e65";
		wait for Clk_period;
		Addr <=  "0001101001011";
		Trees_din <= x"005a0e65";
		wait for Clk_period;
		Addr <=  "0001101001100";
		Trees_din <= x"52feec08";
		wait for Clk_period;
		Addr <=  "0001101001101";
		Trees_din <= x"afffaa04";
		wait for Clk_period;
		Addr <=  "0001101001110";
		Trees_din <= x"00bf0e65";
		wait for Clk_period;
		Addr <=  "0001101001111";
		Trees_din <= x"ff7a0e65";
		wait for Clk_period;
		Addr <=  "0001101010000";
		Trees_din <= x"b9fe0304";
		wait for Clk_period;
		Addr <=  "0001101010001";
		Trees_din <= x"ff860e65";
		wait for Clk_period;
		Addr <=  "0001101010010";
		Trees_din <= x"00ab0e65";
		wait for Clk_period;
		Addr <=  "0001101010011";
		Trees_din <= x"24ff8508";
		wait for Clk_period;
		Addr <=  "0001101010100";
		Trees_din <= x"e7ff3604";
		wait for Clk_period;
		Addr <=  "0001101010101";
		Trees_din <= x"00480e65";
		wait for Clk_period;
		Addr <=  "0001101010110";
		Trees_din <= x"ff2c0e65";
		wait for Clk_period;
		Addr <=  "0001101010111";
		Trees_din <= x"f2029408";
		wait for Clk_period;
		Addr <=  "0001101011000";
		Trees_din <= x"56ff3304";
		wait for Clk_period;
		Addr <=  "0001101011001";
		Trees_din <= x"ffe90e65";
		wait for Clk_period;
		Addr <=  "0001101011010";
		Trees_din <= x"00d50e65";
		wait for Clk_period;
		Addr <=  "0001101011011";
		Trees_din <= x"43ff3d04";
		wait for Clk_period;
		Addr <=  "0001101011100";
		Trees_din <= x"ff590e65";
		wait for Clk_period;
		Addr <=  "0001101011101";
		Trees_din <= x"00790e65";
		wait for Clk_period;
		Addr <=  "0001101011110";
		Trees_din <= x"1dff5040";
		wait for Clk_period;
		Addr <=  "0001101011111";
		Trees_din <= x"7d004520";
		wait for Clk_period;
		Addr <=  "0001101100000";
		Trees_din <= x"c4fef110";
		wait for Clk_period;
		Addr <=  "0001101100001";
		Trees_din <= x"a7ff8508";
		wait for Clk_period;
		Addr <=  "0001101100010";
		Trees_din <= x"71ffc304";
		wait for Clk_period;
		Addr <=  "0001101100011";
		Trees_din <= x"00480e65";
		wait for Clk_period;
		Addr <=  "0001101100100";
		Trees_din <= x"ff7d0e65";
		wait for Clk_period;
		Addr <=  "0001101100101";
		Trees_din <= x"a0fead04";
		wait for Clk_period;
		Addr <=  "0001101100110";
		Trees_din <= x"00090e65";
		wait for Clk_period;
		Addr <=  "0001101100111";
		Trees_din <= x"ff810e65";
		wait for Clk_period;
		Addr <=  "0001101101000";
		Trees_din <= x"cc002f08";
		wait for Clk_period;
		Addr <=  "0001101101001";
		Trees_din <= x"63ffa904";
		wait for Clk_period;
		Addr <=  "0001101101010";
		Trees_din <= x"00700e65";
		wait for Clk_period;
		Addr <=  "0001101101011";
		Trees_din <= x"00230e65";
		wait for Clk_period;
		Addr <=  "0001101101100";
		Trees_din <= x"c9ff9504";
		wait for Clk_period;
		Addr <=  "0001101101101";
		Trees_din <= x"00590e65";
		wait for Clk_period;
		Addr <=  "0001101101110";
		Trees_din <= x"ffbf0e65";
		wait for Clk_period;
		Addr <=  "0001101101111";
		Trees_din <= x"65ff6610";
		wait for Clk_period;
		Addr <=  "0001101110000";
		Trees_din <= x"45fe2a08";
		wait for Clk_period;
		Addr <=  "0001101110001";
		Trees_din <= x"a4ff2704";
		wait for Clk_period;
		Addr <=  "0001101110010";
		Trees_din <= x"00af0e65";
		wait for Clk_period;
		Addr <=  "0001101110011";
		Trees_din <= x"ffaa0e65";
		wait for Clk_period;
		Addr <=  "0001101110100";
		Trees_din <= x"7afee404";
		wait for Clk_period;
		Addr <=  "0001101110101";
		Trees_din <= x"00210e65";
		wait for Clk_period;
		Addr <=  "0001101110110";
		Trees_din <= x"ff380e65";
		wait for Clk_period;
		Addr <=  "0001101110111";
		Trees_din <= x"dfff6508";
		wait for Clk_period;
		Addr <=  "0001101111000";
		Trees_din <= x"77fee104";
		wait for Clk_period;
		Addr <=  "0001101111001";
		Trees_din <= x"00290e65";
		wait for Clk_period;
		Addr <=  "0001101111010";
		Trees_din <= x"ff560e65";
		wait for Clk_period;
		Addr <=  "0001101111011";
		Trees_din <= x"18ff9904";
		wait for Clk_period;
		Addr <=  "0001101111100";
		Trees_din <= x"00db0e65";
		wait for Clk_period;
		Addr <=  "0001101111101";
		Trees_din <= x"ff9c0e65";
		wait for Clk_period;
		Addr <=  "0001101111110";
		Trees_din <= x"3afee318";
		wait for Clk_period;
		Addr <=  "0001101111111";
		Trees_din <= x"2100130c";
		wait for Clk_period;
		Addr <=  "0001110000000";
		Trees_din <= x"98fdf204";
		wait for Clk_period;
		Addr <=  "0001110000001";
		Trees_din <= x"00790e65";
		wait for Clk_period;
		Addr <=  "0001110000010";
		Trees_din <= x"44ff0204";
		wait for Clk_period;
		Addr <=  "0001110000011";
		Trees_din <= x"002b0e65";
		wait for Clk_period;
		Addr <=  "0001110000100";
		Trees_din <= x"ff480e65";
		wait for Clk_period;
		Addr <=  "0001110000101";
		Trees_din <= x"26008b08";
		wait for Clk_period;
		Addr <=  "0001110000110";
		Trees_din <= x"b6ff5104";
		wait for Clk_period;
		Addr <=  "0001110000111";
		Trees_din <= x"00be0e65";
		wait for Clk_period;
		Addr <=  "0001110001000";
		Trees_din <= x"00210e65";
		wait for Clk_period;
		Addr <=  "0001110001001";
		Trees_din <= x"ff7a0e65";
		wait for Clk_period;
		Addr <=  "0001110001010";
		Trees_din <= x"9bff2110";
		wait for Clk_period;
		Addr <=  "0001110001011";
		Trees_din <= x"4fff6108";
		wait for Clk_period;
		Addr <=  "0001110001100";
		Trees_din <= x"a9ff8304";
		wait for Clk_period;
		Addr <=  "0001110001101";
		Trees_din <= x"ff960e65";
		wait for Clk_period;
		Addr <=  "0001110001110";
		Trees_din <= x"00750e65";
		wait for Clk_period;
		Addr <=  "0001110001111";
		Trees_din <= x"7ffea904";
		wait for Clk_period;
		Addr <=  "0001110010000";
		Trees_din <= x"00460e65";
		wait for Clk_period;
		Addr <=  "0001110010001";
		Trees_din <= x"ff4e0e65";
		wait for Clk_period;
		Addr <=  "0001110010010";
		Trees_din <= x"6d002608";
		wait for Clk_period;
		Addr <=  "0001110010011";
		Trees_din <= x"29ff3104";
		wait for Clk_period;
		Addr <=  "0001110010100";
		Trees_din <= x"ffbe0e65";
		wait for Clk_period;
		Addr <=  "0001110010101";
		Trees_din <= x"00910e65";
		wait for Clk_period;
		Addr <=  "0001110010110";
		Trees_din <= x"6cff9c04";
		wait for Clk_period;
		Addr <=  "0001110010111";
		Trees_din <= x"ff900e65";
		wait for Clk_period;
		Addr <=  "0001110011000";
		Trees_din <= x"00460e65";
		wait for Clk_period;
		Addr <=  "0001110011001";
		Trees_din <= x"0dff9e78";
		wait for Clk_period;
		Addr <=  "0001110011010";
		Trees_din <= x"24ff8638";
		wait for Clk_period;
		Addr <=  "0001110011011";
		Trees_din <= x"d5fffe18";
		wait for Clk_period;
		Addr <=  "0001110011100";
		Trees_din <= x"86ffc810";
		wait for Clk_period;
		Addr <=  "0001110011101";
		Trees_din <= x"43ff3d08";
		wait for Clk_period;
		Addr <=  "0001110011110";
		Trees_din <= x"cbffdb04";
		wait for Clk_period;
		Addr <=  "0001110011111";
		Trees_din <= x"ffa51021";
		wait for Clk_period;
		Addr <=  "0001110100000";
		Trees_din <= x"003d1021";
		wait for Clk_period;
		Addr <=  "0001110100001";
		Trees_din <= x"b3ff4304";
		wait for Clk_period;
		Addr <=  "0001110100010";
		Trees_din <= x"00091021";
		wait for Clk_period;
		Addr <=  "0001110100011";
		Trees_din <= x"00871021";
		wait for Clk_period;
		Addr <=  "0001110100100";
		Trees_din <= x"65ffeb04";
		wait for Clk_period;
		Addr <=  "0001110100101";
		Trees_din <= x"ff4f1021";
		wait for Clk_period;
		Addr <=  "0001110100110";
		Trees_din <= x"00521021";
		wait for Clk_period;
		Addr <=  "0001110100111";
		Trees_din <= x"0bffe510";
		wait for Clk_period;
		Addr <=  "0001110101000";
		Trees_din <= x"69ff1408";
		wait for Clk_period;
		Addr <=  "0001110101001";
		Trees_din <= x"5eff9304";
		wait for Clk_period;
		Addr <=  "0001110101010";
		Trees_din <= x"fff71021";
		wait for Clk_period;
		Addr <=  "0001110101011";
		Trees_din <= x"ff2c1021";
		wait for Clk_period;
		Addr <=  "0001110101100";
		Trees_din <= x"d2fedd04";
		wait for Clk_period;
		Addr <=  "0001110101101";
		Trees_din <= x"003c1021";
		wait for Clk_period;
		Addr <=  "0001110101110";
		Trees_din <= x"ffbe1021";
		wait for Clk_period;
		Addr <=  "0001110101111";
		Trees_din <= x"e0ffb908";
		wait for Clk_period;
		Addr <=  "0001110110000";
		Trees_din <= x"33fffd04";
		wait for Clk_period;
		Addr <=  "0001110110001";
		Trees_din <= x"ff511021";
		wait for Clk_period;
		Addr <=  "0001110110010";
		Trees_din <= x"00641021";
		wait for Clk_period;
		Addr <=  "0001110110011";
		Trees_din <= x"c3ffec04";
		wait for Clk_period;
		Addr <=  "0001110110100";
		Trees_din <= x"ff6e1021";
		wait for Clk_period;
		Addr <=  "0001110110101";
		Trees_din <= x"008e1021";
		wait for Clk_period;
		Addr <=  "0001110110110";
		Trees_din <= x"1aff1920";
		wait for Clk_period;
		Addr <=  "0001110110111";
		Trees_din <= x"d8003e10";
		wait for Clk_period;
		Addr <=  "0001110111000";
		Trees_din <= x"5fff0008";
		wait for Clk_period;
		Addr <=  "0001110111001";
		Trees_din <= x"80ff7704";
		wait for Clk_period;
		Addr <=  "0001110111010";
		Trees_din <= x"00281021";
		wait for Clk_period;
		Addr <=  "0001110111011";
		Trees_din <= x"ff9f1021";
		wait for Clk_period;
		Addr <=  "0001110111100";
		Trees_din <= x"cafda104";
		wait for Clk_period;
		Addr <=  "0001110111101";
		Trees_din <= x"ff8a1021";
		wait for Clk_period;
		Addr <=  "0001110111110";
		Trees_din <= x"005d1021";
		wait for Clk_period;
		Addr <=  "0001110111111";
		Trees_din <= x"b3ff5108";
		wait for Clk_period;
		Addr <=  "0001111000000";
		Trees_din <= x"40004504";
		wait for Clk_period;
		Addr <=  "0001111000001";
		Trees_din <= x"ffe31021";
		wait for Clk_period;
		Addr <=  "0001111000010";
		Trees_din <= x"ff6d1021";
		wait for Clk_period;
		Addr <=  "0001111000011";
		Trees_din <= x"49fff804";
		wait for Clk_period;
		Addr <=  "0001111000100";
		Trees_din <= x"fff21021";
		wait for Clk_period;
		Addr <=  "0001111000101";
		Trees_din <= x"00711021";
		wait for Clk_period;
		Addr <=  "0001111000110";
		Trees_din <= x"32fee210";
		wait for Clk_period;
		Addr <=  "0001111000111";
		Trees_din <= x"28fe8508";
		wait for Clk_period;
		Addr <=  "0001111001000";
		Trees_din <= x"65ff6f04";
		wait for Clk_period;
		Addr <=  "0001111001001";
		Trees_din <= x"ff4e1021";
		wait for Clk_period;
		Addr <=  "0001111001010";
		Trees_din <= x"fffb1021";
		wait for Clk_period;
		Addr <=  "0001111001011";
		Trees_din <= x"27008704";
		wait for Clk_period;
		Addr <=  "0001111001100";
		Trees_din <= x"00a81021";
		wait for Clk_period;
		Addr <=  "0001111001101";
		Trees_din <= x"ff711021";
		wait for Clk_period;
		Addr <=  "0001111001110";
		Trees_din <= x"f9fec708";
		wait for Clk_period;
		Addr <=  "0001111001111";
		Trees_din <= x"6effec04";
		wait for Clk_period;
		Addr <=  "0001111010000";
		Trees_din <= x"008a1021";
		wait for Clk_period;
		Addr <=  "0001111010001";
		Trees_din <= x"ff721021";
		wait for Clk_period;
		Addr <=  "0001111010010";
		Trees_din <= x"05009504";
		wait for Clk_period;
		Addr <=  "0001111010011";
		Trees_din <= x"004b1021";
		wait for Clk_period;
		Addr <=  "0001111010100";
		Trees_din <= x"ff9d1021";
		wait for Clk_period;
		Addr <=  "0001111010101";
		Trees_din <= x"5dffee40";
		wait for Clk_period;
		Addr <=  "0001111010110";
		Trees_din <= x"d9ffd320";
		wait for Clk_period;
		Addr <=  "0001111010111";
		Trees_din <= x"8900c510";
		wait for Clk_period;
		Addr <=  "0001111011000";
		Trees_din <= x"1dff5008";
		wait for Clk_period;
		Addr <=  "0001111011001";
		Trees_din <= x"24ff0304";
		wait for Clk_period;
		Addr <=  "0001111011010";
		Trees_din <= x"ff9d1021";
		wait for Clk_period;
		Addr <=  "0001111011011";
		Trees_din <= x"00651021";
		wait for Clk_period;
		Addr <=  "0001111011100";
		Trees_din <= x"91ffcc04";
		wait for Clk_period;
		Addr <=  "0001111011101";
		Trees_din <= x"ffbf1021";
		wait for Clk_period;
		Addr <=  "0001111011110";
		Trees_din <= x"00761021";
		wait for Clk_period;
		Addr <=  "0001111011111";
		Trees_din <= x"7a001208";
		wait for Clk_period;
		Addr <=  "0001111100000";
		Trees_din <= x"d3ff3f04";
		wait for Clk_period;
		Addr <=  "0001111100001";
		Trees_din <= x"ff321021";
		wait for Clk_period;
		Addr <=  "0001111100010";
		Trees_din <= x"006c1021";
		wait for Clk_period;
		Addr <=  "0001111100011";
		Trees_din <= x"0efe6b04";
		wait for Clk_period;
		Addr <=  "0001111100100";
		Trees_din <= x"00af1021";
		wait for Clk_period;
		Addr <=  "0001111100101";
		Trees_din <= x"002a1021";
		wait for Clk_period;
		Addr <=  "0001111100110";
		Trees_din <= x"1bffa810";
		wait for Clk_period;
		Addr <=  "0001111100111";
		Trees_din <= x"6e001b08";
		wait for Clk_period;
		Addr <=  "0001111101000";
		Trees_din <= x"20ff7304";
		wait for Clk_period;
		Addr <=  "0001111101001";
		Trees_din <= x"00421021";
		wait for Clk_period;
		Addr <=  "0001111101010";
		Trees_din <= x"ff951021";
		wait for Clk_period;
		Addr <=  "0001111101011";
		Trees_din <= x"6e00b404";
		wait for Clk_period;
		Addr <=  "0001111101100";
		Trees_din <= x"008c1021";
		wait for Clk_period;
		Addr <=  "0001111101101";
		Trees_din <= x"ffcc1021";
		wait for Clk_period;
		Addr <=  "0001111101110";
		Trees_din <= x"efffcd08";
		wait for Clk_period;
		Addr <=  "0001111101111";
		Trees_din <= x"2a004c04";
		wait for Clk_period;
		Addr <=  "0001111110000";
		Trees_din <= x"00231021";
		wait for Clk_period;
		Addr <=  "0001111110001";
		Trees_din <= x"ff611021";
		wait for Clk_period;
		Addr <=  "0001111110010";
		Trees_din <= x"7bffcd04";
		wait for Clk_period;
		Addr <=  "0001111110011";
		Trees_din <= x"ff271021";
		wait for Clk_period;
		Addr <=  "0001111110100";
		Trees_din <= x"005d1021";
		wait for Clk_period;
		Addr <=  "0001111110101";
		Trees_din <= x"d5009d20";
		wait for Clk_period;
		Addr <=  "0001111110110";
		Trees_din <= x"1fffe810";
		wait for Clk_period;
		Addr <=  "0001111110111";
		Trees_din <= x"d2ff7808";
		wait for Clk_period;
		Addr <=  "0001111111000";
		Trees_din <= x"81ff4504";
		wait for Clk_period;
		Addr <=  "0001111111001";
		Trees_din <= x"00291021";
		wait for Clk_period;
		Addr <=  "0001111111010";
		Trees_din <= x"00951021";
		wait for Clk_period;
		Addr <=  "0001111111011";
		Trees_din <= x"bbff9704";
		wait for Clk_period;
		Addr <=  "0001111111100";
		Trees_din <= x"004c1021";
		wait for Clk_period;
		Addr <=  "0001111111101";
		Trees_din <= x"ff171021";
		wait for Clk_period;
		Addr <=  "0001111111110";
		Trees_din <= x"03ffb508";
		wait for Clk_period;
		Addr <=  "0001111111111";
		Trees_din <= x"6cff6704";
		wait for Clk_period;
		Addr <=  "0010000000000";
		Trees_din <= x"ffab1021";
		wait for Clk_period;
		Addr <=  "0010000000001";
		Trees_din <= x"00901021";
		wait for Clk_period;
		Addr <=  "0010000000010";
		Trees_din <= x"d0009304";
		wait for Clk_period;
		Addr <=  "0010000000011";
		Trees_din <= x"004d1021";
		wait for Clk_period;
		Addr <=  "0010000000100";
		Trees_din <= x"ff7d1021";
		wait for Clk_period;
		Addr <=  "0010000000101";
		Trees_din <= x"1fff7404";
		wait for Clk_period;
		Addr <=  "0010000000110";
		Trees_din <= x"ff4e1021";
		wait for Clk_period;
		Addr <=  "0010000000111";
		Trees_din <= x"ffe41021";
		wait for Clk_period;
		Addr <=  "0010000001000";
		Trees_din <= x"7d004578";
		wait for Clk_period;
		Addr <=  "0010000001001";
		Trees_din <= x"6d005b3c";
		wait for Clk_period;
		Addr <=  "0010000001010";
		Trees_din <= x"dc003c20";
		wait for Clk_period;
		Addr <=  "0010000001011";
		Trees_din <= x"bcff5a10";
		wait for Clk_period;
		Addr <=  "0010000001100";
		Trees_din <= x"74003908";
		wait for Clk_period;
		Addr <=  "0010000001101";
		Trees_din <= x"8ffdf704";
		wait for Clk_period;
		Addr <=  "0010000001110";
		Trees_din <= x"009911ad";
		wait for Clk_period;
		Addr <=  "0010000001111";
		Trees_din <= x"000f11ad";
		wait for Clk_period;
		Addr <=  "0010000010000";
		Trees_din <= x"a5ff8d04";
		wait for Clk_period;
		Addr <=  "0010000010001";
		Trees_din <= x"007111ad";
		wait for Clk_period;
		Addr <=  "0010000010010";
		Trees_din <= x"ff9711ad";
		wait for Clk_period;
		Addr <=  "0010000010011";
		Trees_din <= x"2e006b08";
		wait for Clk_period;
		Addr <=  "0010000010100";
		Trees_din <= x"b3ff9b04";
		wait for Clk_period;
		Addr <=  "0010000010101";
		Trees_din <= x"006211ad";
		wait for Clk_period;
		Addr <=  "0010000010110";
		Trees_din <= x"ffe811ad";
		wait for Clk_period;
		Addr <=  "0010000010111";
		Trees_din <= x"05002604";
		wait for Clk_period;
		Addr <=  "0010000011000";
		Trees_din <= x"ff4311ad";
		wait for Clk_period;
		Addr <=  "0010000011001";
		Trees_din <= x"003511ad";
		wait for Clk_period;
		Addr <=  "0010000011010";
		Trees_din <= x"d7ffe50c";
		wait for Clk_period;
		Addr <=  "0010000011011";
		Trees_din <= x"13002b04";
		wait for Clk_period;
		Addr <=  "0010000011100";
		Trees_din <= x"ffbc11ad";
		wait for Clk_period;
		Addr <=  "0010000011101";
		Trees_din <= x"53ffdb04";
		wait for Clk_period;
		Addr <=  "0010000011110";
		Trees_din <= x"00c211ad";
		wait for Clk_period;
		Addr <=  "0010000011111";
		Trees_din <= x"001e11ad";
		wait for Clk_period;
		Addr <=  "0010000100000";
		Trees_din <= x"aeff4f08";
		wait for Clk_period;
		Addr <=  "0010000100001";
		Trees_din <= x"1dfee604";
		wait for Clk_period;
		Addr <=  "0010000100010";
		Trees_din <= x"001011ad";
		wait for Clk_period;
		Addr <=  "0010000100011";
		Trees_din <= x"ffaf11ad";
		wait for Clk_period;
		Addr <=  "0010000100100";
		Trees_din <= x"97fe9404";
		wait for Clk_period;
		Addr <=  "0010000100101";
		Trees_din <= x"ff7a11ad";
		wait for Clk_period;
		Addr <=  "0010000100110";
		Trees_din <= x"006111ad";
		wait for Clk_period;
		Addr <=  "0010000100111";
		Trees_din <= x"ee003b1c";
		wait for Clk_period;
		Addr <=  "0010000101000";
		Trees_din <= x"f5007e10";
		wait for Clk_period;
		Addr <=  "0010000101001";
		Trees_din <= x"f6ffbd08";
		wait for Clk_period;
		Addr <=  "0010000101010";
		Trees_din <= x"76000004";
		wait for Clk_period;
		Addr <=  "0010000101011";
		Trees_din <= x"ffdb11ad";
		wait for Clk_period;
		Addr <=  "0010000101100";
		Trees_din <= x"ff7911ad";
		wait for Clk_period;
		Addr <=  "0010000101101";
		Trees_din <= x"5dffe104";
		wait for Clk_period;
		Addr <=  "0010000101110";
		Trees_din <= x"00be11ad";
		wait for Clk_period;
		Addr <=  "0010000101111";
		Trees_din <= x"ffd111ad";
		wait for Clk_period;
		Addr <=  "0010000110000";
		Trees_din <= x"86ffa208";
		wait for Clk_period;
		Addr <=  "0010000110001";
		Trees_din <= x"80ffc004";
		wait for Clk_period;
		Addr <=  "0010000110010";
		Trees_din <= x"00cc11ad";
		wait for Clk_period;
		Addr <=  "0010000110011";
		Trees_din <= x"ffdd11ad";
		wait for Clk_period;
		Addr <=  "0010000110100";
		Trees_din <= x"ff7511ad";
		wait for Clk_period;
		Addr <=  "0010000110101";
		Trees_din <= x"20ff3f10";
		wait for Clk_period;
		Addr <=  "0010000110110";
		Trees_din <= x"4ffff008";
		wait for Clk_period;
		Addr <=  "0010000110111";
		Trees_din <= x"87ff1304";
		wait for Clk_period;
		Addr <=  "0010000111000";
		Trees_din <= x"ffd711ad";
		wait for Clk_period;
		Addr <=  "0010000111001";
		Trees_din <= x"00c411ad";
		wait for Clk_period;
		Addr <=  "0010000111010";
		Trees_din <= x"61ff2704";
		wait for Clk_period;
		Addr <=  "0010000111011";
		Trees_din <= x"ff6d11ad";
		wait for Clk_period;
		Addr <=  "0010000111100";
		Trees_din <= x"007711ad";
		wait for Clk_period;
		Addr <=  "0010000111101";
		Trees_din <= x"7dffc308";
		wait for Clk_period;
		Addr <=  "0010000111110";
		Trees_din <= x"cafe9304";
		wait for Clk_period;
		Addr <=  "0010000111111";
		Trees_din <= x"008411ad";
		wait for Clk_period;
		Addr <=  "0010001000000";
		Trees_din <= x"ffe411ad";
		wait for Clk_period;
		Addr <=  "0010001000001";
		Trees_din <= x"54009704";
		wait for Clk_period;
		Addr <=  "0010001000010";
		Trees_din <= x"ff7111ad";
		wait for Clk_period;
		Addr <=  "0010001000011";
		Trees_din <= x"003b11ad";
		wait for Clk_period;
		Addr <=  "0010001000100";
		Trees_din <= x"04ffdd14";
		wait for Clk_period;
		Addr <=  "0010001000101";
		Trees_din <= x"12ffb608";
		wait for Clk_period;
		Addr <=  "0010001000110";
		Trees_din <= x"7affc504";
		wait for Clk_period;
		Addr <=  "0010001000111";
		Trees_din <= x"00bd11ad";
		wait for Clk_period;
		Addr <=  "0010001001000";
		Trees_din <= x"001211ad";
		wait for Clk_period;
		Addr <=  "0010001001001";
		Trees_din <= x"51003c08";
		wait for Clk_period;
		Addr <=  "0010001001010";
		Trees_din <= x"d3ff1404";
		wait for Clk_period;
		Addr <=  "0010001001011";
		Trees_din <= x"ff5c11ad";
		wait for Clk_period;
		Addr <=  "0010001001100";
		Trees_din <= x"002511ad";
		wait for Clk_period;
		Addr <=  "0010001001101";
		Trees_din <= x"009011ad";
		wait for Clk_period;
		Addr <=  "0010001001110";
		Trees_din <= x"91ffdd20";
		wait for Clk_period;
		Addr <=  "0010001001111";
		Trees_din <= x"08fffc10";
		wait for Clk_period;
		Addr <=  "0010001010000";
		Trees_din <= x"bdffc508";
		wait for Clk_period;
		Addr <=  "0010001010001";
		Trees_din <= x"0d002d04";
		wait for Clk_period;
		Addr <=  "0010001010010";
		Trees_din <= x"ff5311ad";
		wait for Clk_period;
		Addr <=  "0010001010011";
		Trees_din <= x"003211ad";
		wait for Clk_period;
		Addr <=  "0010001010100";
		Trees_din <= x"17ffd504";
		wait for Clk_period;
		Addr <=  "0010001010101";
		Trees_din <= x"ffb511ad";
		wait for Clk_period;
		Addr <=  "0010001010110";
		Trees_din <= x"00c111ad";
		wait for Clk_period;
		Addr <=  "0010001010111";
		Trees_din <= x"b6fe9b08";
		wait for Clk_period;
		Addr <=  "0010001011000";
		Trees_din <= x"0bffa304";
		wait for Clk_period;
		Addr <=  "0010001011001";
		Trees_din <= x"00b811ad";
		wait for Clk_period;
		Addr <=  "0010001011010";
		Trees_din <= x"ffe911ad";
		wait for Clk_period;
		Addr <=  "0010001011011";
		Trees_din <= x"03ff5c04";
		wait for Clk_period;
		Addr <=  "0010001011100";
		Trees_din <= x"ff4511ad";
		wait for Clk_period;
		Addr <=  "0010001011101";
		Trees_din <= x"ffa811ad";
		wait for Clk_period;
		Addr <=  "0010001011110";
		Trees_din <= x"9cff7310";
		wait for Clk_period;
		Addr <=  "0010001011111";
		Trees_din <= x"97feb008";
		wait for Clk_period;
		Addr <=  "0010001100000";
		Trees_din <= x"24ff4b04";
		wait for Clk_period;
		Addr <=  "0010001100001";
		Trees_din <= x"fffd11ad";
		wait for Clk_period;
		Addr <=  "0010001100010";
		Trees_din <= x"ff8111ad";
		wait for Clk_period;
		Addr <=  "0010001100011";
		Trees_din <= x"e0ff7104";
		wait for Clk_period;
		Addr <=  "0010001100100";
		Trees_din <= x"00dc11ad";
		wait for Clk_period;
		Addr <=  "0010001100101";
		Trees_din <= x"002a11ad";
		wait for Clk_period;
		Addr <=  "0010001100110";
		Trees_din <= x"4cfe5a04";
		wait for Clk_period;
		Addr <=  "0010001100111";
		Trees_din <= x"008811ad";
		wait for Clk_period;
		Addr <=  "0010001101000";
		Trees_din <= x"d0ffda04";
		wait for Clk_period;
		Addr <=  "0010001101001";
		Trees_din <= x"001511ad";
		wait for Clk_period;
		Addr <=  "0010001101010";
		Trees_din <= x"ff4b11ad";
		wait for Clk_period;
		Addr <=  "0010001101011";
		Trees_din <= x"1efef23c";
		wait for Clk_period;
		Addr <=  "0010001101100";
		Trees_din <= x"2b00a830";
		wait for Clk_period;
		Addr <=  "0010001101101";
		Trees_din <= x"b4ff701c";
		wait for Clk_period;
		Addr <=  "0010001101110";
		Trees_din <= x"91ffee0c";
		wait for Clk_period;
		Addr <=  "0010001101111";
		Trees_din <= x"05ffb904";
		wait for Clk_period;
		Addr <=  "0010001110000";
		Trees_din <= x"00521321";
		wait for Clk_period;
		Addr <=  "0010001110001";
		Trees_din <= x"ddfe4004";
		wait for Clk_period;
		Addr <=  "0010001110010";
		Trees_din <= x"001e1321";
		wait for Clk_period;
		Addr <=  "0010001110011";
		Trees_din <= x"ff531321";
		wait for Clk_period;
		Addr <=  "0010001110100";
		Trees_din <= x"27000408";
		wait for Clk_period;
		Addr <=  "0010001110101";
		Trees_din <= x"75004f04";
		wait for Clk_period;
		Addr <=  "0010001110110";
		Trees_din <= x"00a91321";
		wait for Clk_period;
		Addr <=  "0010001110111";
		Trees_din <= x"00241321";
		wait for Clk_period;
		Addr <=  "0010001111000";
		Trees_din <= x"92fe9904";
		wait for Clk_period;
		Addr <=  "0010001111001";
		Trees_din <= x"002e1321";
		wait for Clk_period;
		Addr <=  "0010001111010";
		Trees_din <= x"ff601321";
		wait for Clk_period;
		Addr <=  "0010001111011";
		Trees_din <= x"84ff9a08";
		wait for Clk_period;
		Addr <=  "0010001111100";
		Trees_din <= x"81ff7e04";
		wait for Clk_period;
		Addr <=  "0010001111101";
		Trees_din <= x"00271321";
		wait for Clk_period;
		Addr <=  "0010001111110";
		Trees_din <= x"00ac1321";
		wait for Clk_period;
		Addr <=  "0010001111111";
		Trees_din <= x"a9ffb904";
		wait for Clk_period;
		Addr <=  "0010010000000";
		Trees_din <= x"ff621321";
		wait for Clk_period;
		Addr <=  "0010010000001";
		Trees_din <= x"75002504";
		wait for Clk_period;
		Addr <=  "0010010000010";
		Trees_din <= x"008c1321";
		wait for Clk_period;
		Addr <=  "0010010000011";
		Trees_din <= x"ffa81321";
		wait for Clk_period;
		Addr <=  "0010010000100";
		Trees_din <= x"b1ff3f08";
		wait for Clk_period;
		Addr <=  "0010010000101";
		Trees_din <= x"42ff5304";
		wait for Clk_period;
		Addr <=  "0010010000110";
		Trees_din <= x"00cc1321";
		wait for Clk_period;
		Addr <=  "0010010000111";
		Trees_din <= x"00311321";
		wait for Clk_period;
		Addr <=  "0010010001000";
		Trees_din <= x"ff8f1321";
		wait for Clk_period;
		Addr <=  "0010010001001";
		Trees_din <= x"2bff8940";
		wait for Clk_period;
		Addr <=  "0010010001010";
		Trees_din <= x"b6ff7220";
		wait for Clk_period;
		Addr <=  "0010010001011";
		Trees_din <= x"9d004f10";
		wait for Clk_period;
		Addr <=  "0010010001100";
		Trees_din <= x"e1005208";
		wait for Clk_period;
		Addr <=  "0010010001101";
		Trees_din <= x"45ff1604";
		wait for Clk_period;
		Addr <=  "0010010001110";
		Trees_din <= x"000a1321";
		wait for Clk_period;
		Addr <=  "0010010001111";
		Trees_din <= x"00541321";
		wait for Clk_period;
		Addr <=  "0010010010000";
		Trees_din <= x"7dff7704";
		wait for Clk_period;
		Addr <=  "0010010010001";
		Trees_din <= x"00331321";
		wait for Clk_period;
		Addr <=  "0010010010010";
		Trees_din <= x"ff7c1321";
		wait for Clk_period;
		Addr <=  "0010010010011";
		Trees_din <= x"61ffe908";
		wait for Clk_period;
		Addr <=  "0010010010100";
		Trees_din <= x"bf001b04";
		wait for Clk_period;
		Addr <=  "0010010010101";
		Trees_din <= x"ff311321";
		wait for Clk_period;
		Addr <=  "0010010010110";
		Trees_din <= x"003b1321";
		wait for Clk_period;
		Addr <=  "0010010010111";
		Trees_din <= x"52ff4404";
		wait for Clk_period;
		Addr <=  "0010010011000";
		Trees_din <= x"fff91321";
		wait for Clk_period;
		Addr <=  "0010010011001";
		Trees_din <= x"00821321";
		wait for Clk_period;
		Addr <=  "0010010011010";
		Trees_din <= x"b2001710";
		wait for Clk_period;
		Addr <=  "0010010011011";
		Trees_din <= x"62ff9308";
		wait for Clk_period;
		Addr <=  "0010010011100";
		Trees_din <= x"cbffd104";
		wait for Clk_period;
		Addr <=  "0010010011101";
		Trees_din <= x"ff7e1321";
		wait for Clk_period;
		Addr <=  "0010010011110";
		Trees_din <= x"ffd61321";
		wait for Clk_period;
		Addr <=  "0010010011111";
		Trees_din <= x"65ff7804";
		wait for Clk_period;
		Addr <=  "0010010100000";
		Trees_din <= x"ffba1321";
		wait for Clk_period;
		Addr <=  "0010010100001";
		Trees_din <= x"00951321";
		wait for Clk_period;
		Addr <=  "0010010100010";
		Trees_din <= x"da002008";
		wait for Clk_period;
		Addr <=  "0010010100011";
		Trees_din <= x"33ff3004";
		wait for Clk_period;
		Addr <=  "0010010100100";
		Trees_din <= x"ffc11321";
		wait for Clk_period;
		Addr <=  "0010010100101";
		Trees_din <= x"00901321";
		wait for Clk_period;
		Addr <=  "0010010100110";
		Trees_din <= x"baff6b04";
		wait for Clk_period;
		Addr <=  "0010010100111";
		Trees_din <= x"008d1321";
		wait for Clk_period;
		Addr <=  "0010010101000";
		Trees_din <= x"ff621321";
		wait for Clk_period;
		Addr <=  "0010010101001";
		Trees_din <= x"49ffa520";
		wait for Clk_period;
		Addr <=  "0010010101010";
		Trees_din <= x"61ff8a10";
		wait for Clk_period;
		Addr <=  "0010010101011";
		Trees_din <= x"37ffe908";
		wait for Clk_period;
		Addr <=  "0010010101100";
		Trees_din <= x"aafff604";
		wait for Clk_period;
		Addr <=  "0010010101101";
		Trees_din <= x"ff9e1321";
		wait for Clk_period;
		Addr <=  "0010010101110";
		Trees_din <= x"003c1321";
		wait for Clk_period;
		Addr <=  "0010010101111";
		Trees_din <= x"18fee504";
		wait for Clk_period;
		Addr <=  "0010010110000";
		Trees_din <= x"ff9d1321";
		wait for Clk_period;
		Addr <=  "0010010110001";
		Trees_din <= x"00751321";
		wait for Clk_period;
		Addr <=  "0010010110010";
		Trees_din <= x"17004508";
		wait for Clk_period;
		Addr <=  "0010010110011";
		Trees_din <= x"a3fef604";
		wait for Clk_period;
		Addr <=  "0010010110100";
		Trees_din <= x"ff751321";
		wait for Clk_period;
		Addr <=  "0010010110101";
		Trees_din <= x"00571321";
		wait for Clk_period;
		Addr <=  "0010010110110";
		Trees_din <= x"e1ff9f04";
		wait for Clk_period;
		Addr <=  "0010010110111";
		Trees_din <= x"00801321";
		wait for Clk_period;
		Addr <=  "0010010111000";
		Trees_din <= x"ff3c1321";
		wait for Clk_period;
		Addr <=  "0010010111001";
		Trees_din <= x"9bfedb10";
		wait for Clk_period;
		Addr <=  "0010010111010";
		Trees_din <= x"d5ff9c08";
		wait for Clk_period;
		Addr <=  "0010010111011";
		Trees_din <= x"1fffeb04";
		wait for Clk_period;
		Addr <=  "0010010111100";
		Trees_din <= x"000f1321";
		wait for Clk_period;
		Addr <=  "0010010111101";
		Trees_din <= x"00d11321";
		wait for Clk_period;
		Addr <=  "0010010111110";
		Trees_din <= x"12ff7904";
		wait for Clk_period;
		Addr <=  "0010010111111";
		Trees_din <= x"00281321";
		wait for Clk_period;
		Addr <=  "0010011000000";
		Trees_din <= x"ffb21321";
		wait for Clk_period;
		Addr <=  "0010011000001";
		Trees_din <= x"5c001308";
		wait for Clk_period;
		Addr <=  "0010011000010";
		Trees_din <= x"95ffaf04";
		wait for Clk_period;
		Addr <=  "0010011000011";
		Trees_din <= x"005c1321";
		wait for Clk_period;
		Addr <=  "0010011000100";
		Trees_din <= x"00091321";
		wait for Clk_period;
		Addr <=  "0010011000101";
		Trees_din <= x"c1fe7a04";
		wait for Clk_period;
		Addr <=  "0010011000110";
		Trees_din <= x"00651321";
		wait for Clk_period;
		Addr <=  "0010011000111";
		Trees_din <= x"000c1321";
		wait for Clk_period;
		Addr <=  "0010011001000";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0010011001001";
		Trees_din <= x"ddfee470";
		wait for Clk_period;
		Addr <=  "0010011001010";
		Trees_din <= x"0dff5030";
		wait for Clk_period;
		Addr <=  "0010011001011";
		Trees_din <= x"7eff1d20";
		wait for Clk_period;
		Addr <=  "0010011001100";
		Trees_din <= x"05fffa10";
		wait for Clk_period;
		Addr <=  "0010011001101";
		Trees_din <= x"36ff4808";
		wait for Clk_period;
		Addr <=  "0010011001110";
		Trees_din <= x"5effa504";
		wait for Clk_period;
		Addr <=  "0010011001111";
		Trees_din <= x"ff4d1501";
		wait for Clk_period;
		Addr <=  "0010011010000";
		Trees_din <= x"002d1501";
		wait for Clk_period;
		Addr <=  "0010011010001";
		Trees_din <= x"8afedc04";
		wait for Clk_period;
		Addr <=  "0010011010010";
		Trees_din <= x"ff841501";
		wait for Clk_period;
		Addr <=  "0010011010011";
		Trees_din <= x"007d1501";
		wait for Clk_period;
		Addr <=  "0010011010100";
		Trees_din <= x"bbfecb08";
		wait for Clk_period;
		Addr <=  "0010011010101";
		Trees_din <= x"4cff4304";
		wait for Clk_period;
		Addr <=  "0010011010110";
		Trees_din <= x"009a1501";
		wait for Clk_period;
		Addr <=  "0010011010111";
		Trees_din <= x"ff711501";
		wait for Clk_period;
		Addr <=  "0010011011000";
		Trees_din <= x"a6ffbf04";
		wait for Clk_period;
		Addr <=  "0010011011001";
		Trees_din <= x"ff621501";
		wait for Clk_period;
		Addr <=  "0010011011010";
		Trees_din <= x"ffd01501";
		wait for Clk_period;
		Addr <=  "0010011011011";
		Trees_din <= x"6effd804";
		wait for Clk_period;
		Addr <=  "0010011011100";
		Trees_din <= x"ff601501";
		wait for Clk_period;
		Addr <=  "0010011011101";
		Trees_din <= x"fdff9e08";
		wait for Clk_period;
		Addr <=  "0010011011110";
		Trees_din <= x"81ffb304";
		wait for Clk_period;
		Addr <=  "0010011011111";
		Trees_din <= x"ffa41501";
		wait for Clk_period;
		Addr <=  "0010011100000";
		Trees_din <= x"00891501";
		wait for Clk_period;
		Addr <=  "0010011100001";
		Trees_din <= x"00bc1501";
		wait for Clk_period;
		Addr <=  "0010011100010";
		Trees_din <= x"27ffd220";
		wait for Clk_period;
		Addr <=  "0010011100011";
		Trees_din <= x"a4ff5010";
		wait for Clk_period;
		Addr <=  "0010011100100";
		Trees_din <= x"b8ff7608";
		wait for Clk_period;
		Addr <=  "0010011100101";
		Trees_din <= x"68ff0b04";
		wait for Clk_period;
		Addr <=  "0010011100110";
		Trees_din <= x"ff441501";
		wait for Clk_period;
		Addr <=  "0010011100111";
		Trees_din <= x"000e1501";
		wait for Clk_period;
		Addr <=  "0010011101000";
		Trees_din <= x"23ffc204";
		wait for Clk_period;
		Addr <=  "0010011101001";
		Trees_din <= x"00711501";
		wait for Clk_period;
		Addr <=  "0010011101010";
		Trees_din <= x"ff7b1501";
		wait for Clk_period;
		Addr <=  "0010011101011";
		Trees_din <= x"a4ffb808";
		wait for Clk_period;
		Addr <=  "0010011101100";
		Trees_din <= x"7d001704";
		wait for Clk_period;
		Addr <=  "0010011101101";
		Trees_din <= x"00881501";
		wait for Clk_period;
		Addr <=  "0010011101110";
		Trees_din <= x"ffcb1501";
		wait for Clk_period;
		Addr <=  "0010011101111";
		Trees_din <= x"1eff8d04";
		wait for Clk_period;
		Addr <=  "0010011110000";
		Trees_din <= x"ff581501";
		wait for Clk_period;
		Addr <=  "0010011110001";
		Trees_din <= x"00411501";
		wait for Clk_period;
		Addr <=  "0010011110010";
		Trees_din <= x"1fff3a10";
		wait for Clk_period;
		Addr <=  "0010011110011";
		Trees_din <= x"dcffea08";
		wait for Clk_period;
		Addr <=  "0010011110100";
		Trees_din <= x"72ffdd04";
		wait for Clk_period;
		Addr <=  "0010011110101";
		Trees_din <= x"ffe31501";
		wait for Clk_period;
		Addr <=  "0010011110110";
		Trees_din <= x"00b01501";
		wait for Clk_period;
		Addr <=  "0010011110111";
		Trees_din <= x"61ff5804";
		wait for Clk_period;
		Addr <=  "0010011111000";
		Trees_din <= x"ff561501";
		wait for Clk_period;
		Addr <=  "0010011111001";
		Trees_din <= x"005a1501";
		wait for Clk_period;
		Addr <=  "0010011111010";
		Trees_din <= x"6effc008";
		wait for Clk_period;
		Addr <=  "0010011111011";
		Trees_din <= x"c3ffb904";
		wait for Clk_period;
		Addr <=  "0010011111100";
		Trees_din <= x"007a1501";
		wait for Clk_period;
		Addr <=  "0010011111101";
		Trees_din <= x"ffda1501";
		wait for Clk_period;
		Addr <=  "0010011111110";
		Trees_din <= x"69ff0d04";
		wait for Clk_period;
		Addr <=  "0010011111111";
		Trees_din <= x"00051501";
		wait for Clk_period;
		Addr <=  "0010100000000";
		Trees_din <= x"ff801501";
		wait for Clk_period;
		Addr <=  "0010100000001";
		Trees_din <= x"65ff5140";
		wait for Clk_period;
		Addr <=  "0010100000010";
		Trees_din <= x"1fff7920";
		wait for Clk_period;
		Addr <=  "0010100000011";
		Trees_din <= x"1bff8310";
		wait for Clk_period;
		Addr <=  "0010100000100";
		Trees_din <= x"9fffda08";
		wait for Clk_period;
		Addr <=  "0010100000101";
		Trees_din <= x"fcff9604";
		wait for Clk_period;
		Addr <=  "0010100000110";
		Trees_din <= x"00961501";
		wait for Clk_period;
		Addr <=  "0010100000111";
		Trees_din <= x"ffcd1501";
		wait for Clk_period;
		Addr <=  "0010100001000";
		Trees_din <= x"f7ff0d04";
		wait for Clk_period;
		Addr <=  "0010100001001";
		Trees_din <= x"00731501";
		wait for Clk_period;
		Addr <=  "0010100001010";
		Trees_din <= x"ff4a1501";
		wait for Clk_period;
		Addr <=  "0010100001011";
		Trees_din <= x"40003908";
		wait for Clk_period;
		Addr <=  "0010100001100";
		Trees_din <= x"7efe8304";
		wait for Clk_period;
		Addr <=  "0010100001101";
		Trees_din <= x"ffb71501";
		wait for Clk_period;
		Addr <=  "0010100001110";
		Trees_din <= x"004f1501";
		wait for Clk_period;
		Addr <=  "0010100001111";
		Trees_din <= x"69ff9404";
		wait for Clk_period;
		Addr <=  "0010100010000";
		Trees_din <= x"ff851501";
		wait for Clk_period;
		Addr <=  "0010100010001";
		Trees_din <= x"00231501";
		wait for Clk_period;
		Addr <=  "0010100010010";
		Trees_din <= x"5bffdb10";
		wait for Clk_period;
		Addr <=  "0010100010011";
		Trees_din <= x"00ff7e08";
		wait for Clk_period;
		Addr <=  "0010100010100";
		Trees_din <= x"6bfe9304";
		wait for Clk_period;
		Addr <=  "0010100010101";
		Trees_din <= x"ffba1501";
		wait for Clk_period;
		Addr <=  "0010100010110";
		Trees_din <= x"001b1501";
		wait for Clk_period;
		Addr <=  "0010100010111";
		Trees_din <= x"a7ff6104";
		wait for Clk_period;
		Addr <=  "0010100011000";
		Trees_din <= x"fff71501";
		wait for Clk_period;
		Addr <=  "0010100011001";
		Trees_din <= x"ff931501";
		wait for Clk_period;
		Addr <=  "0010100011010";
		Trees_din <= x"01fe9c08";
		wait for Clk_period;
		Addr <=  "0010100011011";
		Trees_din <= x"80ff6004";
		wait for Clk_period;
		Addr <=  "0010100011100";
		Trees_din <= x"00761501";
		wait for Clk_period;
		Addr <=  "0010100011101";
		Trees_din <= x"ff691501";
		wait for Clk_period;
		Addr <=  "0010100011110";
		Trees_din <= x"33ffed04";
		wait for Clk_period;
		Addr <=  "0010100011111";
		Trees_din <= x"00c01501";
		wait for Clk_period;
		Addr <=  "0010100100000";
		Trees_din <= x"ff861501";
		wait for Clk_period;
		Addr <=  "0010100100001";
		Trees_din <= x"1f005520";
		wait for Clk_period;
		Addr <=  "0010100100010";
		Trees_din <= x"3dfff410";
		wait for Clk_period;
		Addr <=  "0010100100011";
		Trees_din <= x"5a004508";
		wait for Clk_period;
		Addr <=  "0010100100100";
		Trees_din <= x"62ff9004";
		wait for Clk_period;
		Addr <=  "0010100100101";
		Trees_din <= x"ffc01501";
		wait for Clk_period;
		Addr <=  "0010100100110";
		Trees_din <= x"00871501";
		wait for Clk_period;
		Addr <=  "0010100100111";
		Trees_din <= x"d1ff9c04";
		wait for Clk_period;
		Addr <=  "0010100101000";
		Trees_din <= x"00431501";
		wait for Clk_period;
		Addr <=  "0010100101001";
		Trees_din <= x"ffb81501";
		wait for Clk_period;
		Addr <=  "0010100101010";
		Trees_din <= x"24ff0d08";
		wait for Clk_period;
		Addr <=  "0010100101011";
		Trees_din <= x"c9ffb904";
		wait for Clk_period;
		Addr <=  "0010100101100";
		Trees_din <= x"00761501";
		wait for Clk_period;
		Addr <=  "0010100101101";
		Trees_din <= x"ff3e1501";
		wait for Clk_period;
		Addr <=  "0010100101110";
		Trees_din <= x"00ffd504";
		wait for Clk_period;
		Addr <=  "0010100101111";
		Trees_din <= x"006c1501";
		wait for Clk_period;
		Addr <=  "0010100110000";
		Trees_din <= x"ffcd1501";
		wait for Clk_period;
		Addr <=  "0010100110001";
		Trees_din <= x"d7008310";
		wait for Clk_period;
		Addr <=  "0010100110010";
		Trees_din <= x"deffe008";
		wait for Clk_period;
		Addr <=  "0010100110011";
		Trees_din <= x"aeff1604";
		wait for Clk_period;
		Addr <=  "0010100110100";
		Trees_din <= x"00281501";
		wait for Clk_period;
		Addr <=  "0010100110101";
		Trees_din <= x"ff541501";
		wait for Clk_period;
		Addr <=  "0010100110110";
		Trees_din <= x"f202d504";
		wait for Clk_period;
		Addr <=  "0010100110111";
		Trees_din <= x"00721501";
		wait for Clk_period;
		Addr <=  "0010100111000";
		Trees_din <= x"ffb81501";
		wait for Clk_period;
		Addr <=  "0010100111001";
		Trees_din <= x"cc004708";
		wait for Clk_period;
		Addr <=  "0010100111010";
		Trees_din <= x"32ff0104";
		wait for Clk_period;
		Addr <=  "0010100111011";
		Trees_din <= x"001a1501";
		wait for Clk_period;
		Addr <=  "0010100111100";
		Trees_din <= x"ff4c1501";
		wait for Clk_period;
		Addr <=  "0010100111101";
		Trees_din <= x"8dfd5b04";
		wait for Clk_period;
		Addr <=  "0010100111110";
		Trees_din <= x"00391501";
		wait for Clk_period;
		Addr <=  "0010100111111";
		Trees_din <= x"ff321501";
		wait for Clk_period;
		Addr <=  "0010101000000";
		Trees_din <= x"c8fff464";
		wait for Clk_period;
		Addr <=  "0010101000001";
		Trees_din <= x"2fffe834";
		wait for Clk_period;
		Addr <=  "0010101000010";
		Trees_din <= x"44005b18";
		wait for Clk_period;
		Addr <=  "0010101000011";
		Trees_din <= x"5aff9308";
		wait for Clk_period;
		Addr <=  "0010101000100";
		Trees_din <= x"d1ff5004";
		wait for Clk_period;
		Addr <=  "0010101000101";
		Trees_din <= x"ff4e16b5";
		wait for Clk_period;
		Addr <=  "0010101000110";
		Trees_din <= x"ffe516b5";
		wait for Clk_period;
		Addr <=  "0010101000111";
		Trees_din <= x"50fed708";
		wait for Clk_period;
		Addr <=  "0010101001000";
		Trees_din <= x"53ff7404";
		wait for Clk_period;
		Addr <=  "0010101001001";
		Trees_din <= x"002316b5";
		wait for Clk_period;
		Addr <=  "0010101001010";
		Trees_din <= x"ff8516b5";
		wait for Clk_period;
		Addr <=  "0010101001011";
		Trees_din <= x"24ff0d04";
		wait for Clk_period;
		Addr <=  "0010101001100";
		Trees_din <= x"ffd816b5";
		wait for Clk_period;
		Addr <=  "0010101001101";
		Trees_din <= x"004016b5";
		wait for Clk_period;
		Addr <=  "0010101001110";
		Trees_din <= x"98fe7a0c";
		wait for Clk_period;
		Addr <=  "0010101001111";
		Trees_din <= x"45ff3f08";
		wait for Clk_period;
		Addr <=  "0010101010000";
		Trees_din <= x"b9fed604";
		wait for Clk_period;
		Addr <=  "0010101010001";
		Trees_din <= x"ffd116b5";
		wait for Clk_period;
		Addr <=  "0010101010010";
		Trees_din <= x"fefd16b5";
		wait for Clk_period;
		Addr <=  "0010101010011";
		Trees_din <= x"005916b5";
		wait for Clk_period;
		Addr <=  "0010101010100";
		Trees_din <= x"b6ffa008";
		wait for Clk_period;
		Addr <=  "0010101010101";
		Trees_din <= x"cafdd604";
		wait for Clk_period;
		Addr <=  "0010101010110";
		Trees_din <= x"ff8b16b5";
		wait for Clk_period;
		Addr <=  "0010101010111";
		Trees_din <= x"004916b5";
		wait for Clk_period;
		Addr <=  "0010101011000";
		Trees_din <= x"4cffbe04";
		wait for Clk_period;
		Addr <=  "0010101011001";
		Trees_din <= x"ff4616b5";
		wait for Clk_period;
		Addr <=  "0010101011010";
		Trees_din <= x"006c16b5";
		wait for Clk_period;
		Addr <=  "0010101011011";
		Trees_din <= x"03ffc81c";
		wait for Clk_period;
		Addr <=  "0010101011100";
		Trees_din <= x"09ff620c";
		wait for Clk_period;
		Addr <=  "0010101011101";
		Trees_din <= x"d9ffac08";
		wait for Clk_period;
		Addr <=  "0010101011110";
		Trees_din <= x"de001d04";
		wait for Clk_period;
		Addr <=  "0010101011111";
		Trees_din <= x"ff9e16b5";
		wait for Clk_period;
		Addr <=  "0010101100000";
		Trees_din <= x"008816b5";
		wait for Clk_period;
		Addr <=  "0010101100001";
		Trees_din <= x"ff4516b5";
		wait for Clk_period;
		Addr <=  "0010101100010";
		Trees_din <= x"afff8108";
		wait for Clk_period;
		Addr <=  "0010101100011";
		Trees_din <= x"d3fee904";
		wait for Clk_period;
		Addr <=  "0010101100100";
		Trees_din <= x"ff7016b5";
		wait for Clk_period;
		Addr <=  "0010101100101";
		Trees_din <= x"005916b5";
		wait for Clk_period;
		Addr <=  "0010101100110";
		Trees_din <= x"beff6e04";
		wait for Clk_period;
		Addr <=  "0010101100111";
		Trees_din <= x"ff9a16b5";
		wait for Clk_period;
		Addr <=  "0010101101000";
		Trees_din <= x"00b016b5";
		wait for Clk_period;
		Addr <=  "0010101101001";
		Trees_din <= x"91feff08";
		wait for Clk_period;
		Addr <=  "0010101101010";
		Trees_din <= x"b5fe8604";
		wait for Clk_period;
		Addr <=  "0010101101011";
		Trees_din <= x"009416b5";
		wait for Clk_period;
		Addr <=  "0010101101100";
		Trees_din <= x"000d16b5";
		wait for Clk_period;
		Addr <=  "0010101101101";
		Trees_din <= x"30ff5104";
		wait for Clk_period;
		Addr <=  "0010101101110";
		Trees_din <= x"002116b5";
		wait for Clk_period;
		Addr <=  "0010101101111";
		Trees_din <= x"4ffee204";
		wait for Clk_period;
		Addr <=  "0010101110000";
		Trees_din <= x"000c16b5";
		wait for Clk_period;
		Addr <=  "0010101110001";
		Trees_din <= x"ff2616b5";
		wait for Clk_period;
		Addr <=  "0010101110010";
		Trees_din <= x"d6004840";
		wait for Clk_period;
		Addr <=  "0010101110011";
		Trees_din <= x"3eff9120";
		wait for Clk_period;
		Addr <=  "0010101110100";
		Trees_din <= x"51ff0710";
		wait for Clk_period;
		Addr <=  "0010101110101";
		Trees_din <= x"75001b08";
		wait for Clk_period;
		Addr <=  "0010101110110";
		Trees_din <= x"49ffcb04";
		wait for Clk_period;
		Addr <=  "0010101110111";
		Trees_din <= x"000316b5";
		wait for Clk_period;
		Addr <=  "0010101111000";
		Trees_din <= x"fefb16b5";
		wait for Clk_period;
		Addr <=  "0010101111001";
		Trees_din <= x"d1ff3c04";
		wait for Clk_period;
		Addr <=  "0010101111010";
		Trees_din <= x"008716b5";
		wait for Clk_period;
		Addr <=  "0010101111011";
		Trees_din <= x"ff9116b5";
		wait for Clk_period;
		Addr <=  "0010101111100";
		Trees_din <= x"99fe6408";
		wait for Clk_period;
		Addr <=  "0010101111101";
		Trees_din <= x"e3fe6b04";
		wait for Clk_period;
		Addr <=  "0010101111110";
		Trees_din <= x"ff5816b5";
		wait for Clk_period;
		Addr <=  "0010101111111";
		Trees_din <= x"000a16b5";
		wait for Clk_period;
		Addr <=  "0010110000000";
		Trees_din <= x"8cffab04";
		wait for Clk_period;
		Addr <=  "0010110000001";
		Trees_din <= x"006516b5";
		wait for Clk_period;
		Addr <=  "0010110000010";
		Trees_din <= x"001e16b5";
		wait for Clk_period;
		Addr <=  "0010110000011";
		Trees_din <= x"9bff3d10";
		wait for Clk_period;
		Addr <=  "0010110000100";
		Trees_din <= x"0fff6a08";
		wait for Clk_period;
		Addr <=  "0010110000101";
		Trees_din <= x"5a003f04";
		wait for Clk_period;
		Addr <=  "0010110000110";
		Trees_din <= x"ff7c16b5";
		wait for Clk_period;
		Addr <=  "0010110000111";
		Trees_din <= x"006d16b5";
		wait for Clk_period;
		Addr <=  "0010110001000";
		Trees_din <= x"afff0604";
		wait for Clk_period;
		Addr <=  "0010110001001";
		Trees_din <= x"007416b5";
		wait for Clk_period;
		Addr <=  "0010110001010";
		Trees_din <= x"ff4e16b5";
		wait for Clk_period;
		Addr <=  "0010110001011";
		Trees_din <= x"5bff8408";
		wait for Clk_period;
		Addr <=  "0010110001100";
		Trees_din <= x"7eff1204";
		wait for Clk_period;
		Addr <=  "0010110001101";
		Trees_din <= x"ffbb16b5";
		wait for Clk_period;
		Addr <=  "0010110001110";
		Trees_din <= x"009416b5";
		wait for Clk_period;
		Addr <=  "0010110001111";
		Trees_din <= x"deffd504";
		wait for Clk_period;
		Addr <=  "0010110010000";
		Trees_din <= x"ff7016b5";
		wait for Clk_period;
		Addr <=  "0010110010001";
		Trees_din <= x"006516b5";
		wait for Clk_period;
		Addr <=  "0010110010010";
		Trees_din <= x"75ff9f1c";
		wait for Clk_period;
		Addr <=  "0010110010011";
		Trees_din <= x"dc004610";
		wait for Clk_period;
		Addr <=  "0010110010100";
		Trees_din <= x"8dff8808";
		wait for Clk_period;
		Addr <=  "0010110010101";
		Trees_din <= x"b5fe6904";
		wait for Clk_period;
		Addr <=  "0010110010110";
		Trees_din <= x"ffbf16b5";
		wait for Clk_period;
		Addr <=  "0010110010111";
		Trees_din <= x"008716b5";
		wait for Clk_period;
		Addr <=  "0010110011000";
		Trees_din <= x"0eff1204";
		wait for Clk_period;
		Addr <=  "0010110011001";
		Trees_din <= x"ffd116b5";
		wait for Clk_period;
		Addr <=  "0010110011010";
		Trees_din <= x"ff3d16b5";
		wait for Clk_period;
		Addr <=  "0010110011011";
		Trees_din <= x"feff7904";
		wait for Clk_period;
		Addr <=  "0010110011100";
		Trees_din <= x"005a16b5";
		wait for Clk_period;
		Addr <=  "0010110011101";
		Trees_din <= x"eeff6604";
		wait for Clk_period;
		Addr <=  "0010110011110";
		Trees_din <= x"ffd016b5";
		wait for Clk_period;
		Addr <=  "0010110011111";
		Trees_din <= x"ff5116b5";
		wait for Clk_period;
		Addr <=  "0010110100000";
		Trees_din <= x"5a013410";
		wait for Clk_period;
		Addr <=  "0010110100001";
		Trees_din <= x"27004708";
		wait for Clk_period;
		Addr <=  "0010110100010";
		Trees_din <= x"90ffcb04";
		wait for Clk_period;
		Addr <=  "0010110100011";
		Trees_din <= x"ffe816b5";
		wait for Clk_period;
		Addr <=  "0010110100100";
		Trees_din <= x"ff8516b5";
		wait for Clk_period;
		Addr <=  "0010110100101";
		Trees_din <= x"3fffdc04";
		wait for Clk_period;
		Addr <=  "0010110100110";
		Trees_din <= x"003616b5";
		wait for Clk_period;
		Addr <=  "0010110100111";
		Trees_din <= x"ff5616b5";
		wait for Clk_period;
		Addr <=  "0010110101000";
		Trees_din <= x"00fee604";
		wait for Clk_period;
		Addr <=  "0010110101001";
		Trees_din <= x"ff6416b5";
		wait for Clk_period;
		Addr <=  "0010110101010";
		Trees_din <= x"b2ff7b04";
		wait for Clk_period;
		Addr <=  "0010110101011";
		Trees_din <= x"ffbf16b5";
		wait for Clk_period;
		Addr <=  "0010110101100";
		Trees_din <= x"00a216b5";
		wait for Clk_period;
		Addr <=  "0010110101101";
		Trees_din <= x"b6ff727c";
		wait for Clk_period;
		Addr <=  "0010110101110";
		Trees_din <= x"1bffb33c";
		wait for Clk_period;
		Addr <=  "0010110101111";
		Trees_din <= x"e0fe5b1c";
		wait for Clk_period;
		Addr <=  "0010110110000";
		Trees_din <= x"ee003a10";
		wait for Clk_period;
		Addr <=  "0010110110001";
		Trees_din <= x"13008108";
		wait for Clk_period;
		Addr <=  "0010110110010";
		Trees_din <= x"2cff8b04";
		wait for Clk_period;
		Addr <=  "0010110110011";
		Trees_din <= x"ff881869";
		wait for Clk_period;
		Addr <=  "0010110110100";
		Trees_din <= x"007b1869";
		wait for Clk_period;
		Addr <=  "0010110110101";
		Trees_din <= x"2bff4c04";
		wait for Clk_period;
		Addr <=  "0010110110110";
		Trees_din <= x"00171869";
		wait for Clk_period;
		Addr <=  "0010110110111";
		Trees_din <= x"ff221869";
		wait for Clk_period;
		Addr <=  "0010110111000";
		Trees_din <= x"a9ff5d04";
		wait for Clk_period;
		Addr <=  "0010110111001";
		Trees_din <= x"00911869";
		wait for Clk_period;
		Addr <=  "0010110111010";
		Trees_din <= x"00ff5f04";
		wait for Clk_period;
		Addr <=  "0010110111011";
		Trees_din <= x"00021869";
		wait for Clk_period;
		Addr <=  "0010110111100";
		Trees_din <= x"ff841869";
		wait for Clk_period;
		Addr <=  "0010110111101";
		Trees_din <= x"63ffe010";
		wait for Clk_period;
		Addr <=  "0010110111110";
		Trees_din <= x"1f005208";
		wait for Clk_period;
		Addr <=  "0010110111111";
		Trees_din <= x"90ff9204";
		wait for Clk_period;
		Addr <=  "0010111000000";
		Trees_din <= x"005d1869";
		wait for Clk_period;
		Addr <=  "0010111000001";
		Trees_din <= x"001d1869";
		wait for Clk_period;
		Addr <=  "0010111000010";
		Trees_din <= x"16feb404";
		wait for Clk_period;
		Addr <=  "0010111000011";
		Trees_din <= x"00591869";
		wait for Clk_period;
		Addr <=  "0010111000100";
		Trees_din <= x"ffd31869";
		wait for Clk_period;
		Addr <=  "0010111000101";
		Trees_din <= x"c4ff2308";
		wait for Clk_period;
		Addr <=  "0010111000110";
		Trees_din <= x"de007804";
		wait for Clk_period;
		Addr <=  "0010111000111";
		Trees_din <= x"ff721869";
		wait for Clk_period;
		Addr <=  "0010111001000";
		Trees_din <= x"00561869";
		wait for Clk_period;
		Addr <=  "0010111001001";
		Trees_din <= x"51ff8404";
		wait for Clk_period;
		Addr <=  "0010111001010";
		Trees_din <= x"ffe51869";
		wait for Clk_period;
		Addr <=  "0010111001011";
		Trees_din <= x"00771869";
		wait for Clk_period;
		Addr <=  "0010111001100";
		Trees_din <= x"06ff5a20";
		wait for Clk_period;
		Addr <=  "0010111001101";
		Trees_din <= x"3cff2610";
		wait for Clk_period;
		Addr <=  "0010111001110";
		Trees_din <= x"5a012508";
		wait for Clk_period;
		Addr <=  "0010111001111";
		Trees_din <= x"32fec304";
		wait for Clk_period;
		Addr <=  "0010111010000";
		Trees_din <= x"ffdb1869";
		wait for Clk_period;
		Addr <=  "0010111010001";
		Trees_din <= x"ff5f1869";
		wait for Clk_period;
		Addr <=  "0010111010010";
		Trees_din <= x"a8ff3504";
		wait for Clk_period;
		Addr <=  "0010111010011";
		Trees_din <= x"ffa51869";
		wait for Clk_period;
		Addr <=  "0010111010100";
		Trees_din <= x"00ac1869";
		wait for Clk_period;
		Addr <=  "0010111010101";
		Trees_din <= x"77ff2708";
		wait for Clk_period;
		Addr <=  "0010111010110";
		Trees_din <= x"e2fe8004";
		wait for Clk_period;
		Addr <=  "0010111010111";
		Trees_din <= x"ff7f1869";
		wait for Clk_period;
		Addr <=  "0010111011000";
		Trees_din <= x"00701869";
		wait for Clk_period;
		Addr <=  "0010111011001";
		Trees_din <= x"b3ff6204";
		wait for Clk_period;
		Addr <=  "0010111011010";
		Trees_din <= x"ff971869";
		wait for Clk_period;
		Addr <=  "0010111011011";
		Trees_din <= x"00561869";
		wait for Clk_period;
		Addr <=  "0010111011100";
		Trees_din <= x"91ff7810";
		wait for Clk_period;
		Addr <=  "0010111011101";
		Trees_din <= x"5bff9f08";
		wait for Clk_period;
		Addr <=  "0010111011110";
		Trees_din <= x"ddfec604";
		wait for Clk_period;
		Addr <=  "0010111011111";
		Trees_din <= x"ff691869";
		wait for Clk_period;
		Addr <=  "0010111100000";
		Trees_din <= x"ffe91869";
		wait for Clk_period;
		Addr <=  "0010111100001";
		Trees_din <= x"9bff3704";
		wait for Clk_period;
		Addr <=  "0010111100010";
		Trees_din <= x"ffe31869";
		wait for Clk_period;
		Addr <=  "0010111100011";
		Trees_din <= x"00811869";
		wait for Clk_period;
		Addr <=  "0010111100100";
		Trees_din <= x"3f003a08";
		wait for Clk_period;
		Addr <=  "0010111100101";
		Trees_din <= x"09ffe904";
		wait for Clk_period;
		Addr <=  "0010111100110";
		Trees_din <= x"006a1869";
		wait for Clk_period;
		Addr <=  "0010111100111";
		Trees_din <= x"000a1869";
		wait for Clk_period;
		Addr <=  "0010111101000";
		Trees_din <= x"57ffb304";
		wait for Clk_period;
		Addr <=  "0010111101001";
		Trees_din <= x"ffd91869";
		wait for Clk_period;
		Addr <=  "0010111101010";
		Trees_din <= x"00861869";
		wait for Clk_period;
		Addr <=  "0010111101011";
		Trees_din <= x"da007b40";
		wait for Clk_period;
		Addr <=  "0010111101100";
		Trees_din <= x"0bfff920";
		wait for Clk_period;
		Addr <=  "0010111101101";
		Trees_din <= x"cbff9a10";
		wait for Clk_period;
		Addr <=  "0010111101110";
		Trees_din <= x"beffb508";
		wait for Clk_period;
		Addr <=  "0010111101111";
		Trees_din <= x"39ff1904";
		wait for Clk_period;
		Addr <=  "0010111110000";
		Trees_din <= x"ff951869";
		wait for Clk_period;
		Addr <=  "0010111110001";
		Trees_din <= x"00761869";
		wait for Clk_period;
		Addr <=  "0010111110010";
		Trees_din <= x"cbff0604";
		wait for Clk_period;
		Addr <=  "0010111110011";
		Trees_din <= x"00751869";
		wait for Clk_period;
		Addr <=  "0010111110100";
		Trees_din <= x"ffc11869";
		wait for Clk_period;
		Addr <=  "0010111110101";
		Trees_din <= x"63ffd608";
		wait for Clk_period;
		Addr <=  "0010111110110";
		Trees_din <= x"d6008104";
		wait for Clk_period;
		Addr <=  "0010111110111";
		Trees_din <= x"00481869";
		wait for Clk_period;
		Addr <=  "0010111111000";
		Trees_din <= x"ffdc1869";
		wait for Clk_period;
		Addr <=  "0010111111001";
		Trees_din <= x"78ff3d04";
		wait for Clk_period;
		Addr <=  "0010111111010";
		Trees_din <= x"ff491869";
		wait for Clk_period;
		Addr <=  "0010111111011";
		Trees_din <= x"00001869";
		wait for Clk_period;
		Addr <=  "0010111111100";
		Trees_din <= x"de008410";
		wait for Clk_period;
		Addr <=  "0010111111101";
		Trees_din <= x"19ff3208";
		wait for Clk_period;
		Addr <=  "0010111111110";
		Trees_din <= x"95ff9104";
		wait for Clk_period;
		Addr <=  "0010111111111";
		Trees_din <= x"ff541869";
		wait for Clk_period;
		Addr <=  "0011000000000";
		Trees_din <= x"ffe51869";
		wait for Clk_period;
		Addr <=  "0011000000001";
		Trees_din <= x"f0ff3004";
		wait for Clk_period;
		Addr <=  "0011000000010";
		Trees_din <= x"ff901869";
		wait for Clk_period;
		Addr <=  "0011000000011";
		Trees_din <= x"000e1869";
		wait for Clk_period;
		Addr <=  "0011000000100";
		Trees_din <= x"7affa908";
		wait for Clk_period;
		Addr <=  "0011000000101";
		Trees_din <= x"f6fe9e04";
		wait for Clk_period;
		Addr <=  "0011000000110";
		Trees_din <= x"ff9f1869";
		wait for Clk_period;
		Addr <=  "0011000000111";
		Trees_din <= x"00ac1869";
		wait for Clk_period;
		Addr <=  "0011000001000";
		Trees_din <= x"12ff6b04";
		wait for Clk_period;
		Addr <=  "0011000001001";
		Trees_din <= x"00671869";
		wait for Clk_period;
		Addr <=  "0011000001010";
		Trees_din <= x"ff701869";
		wait for Clk_period;
		Addr <=  "0011000001011";
		Trees_din <= x"75ffff14";
		wait for Clk_period;
		Addr <=  "0011000001100";
		Trees_din <= x"04004a0c";
		wait for Clk_period;
		Addr <=  "0011000001101";
		Trees_din <= x"4afede04";
		wait for Clk_period;
		Addr <=  "0011000001110";
		Trees_din <= x"ff8e1869";
		wait for Clk_period;
		Addr <=  "0011000001111";
		Trees_din <= x"28ff0904";
		wait for Clk_period;
		Addr <=  "0011000010000";
		Trees_din <= x"fff91869";
		wait for Clk_period;
		Addr <=  "0011000010001";
		Trees_din <= x"009a1869";
		wait for Clk_period;
		Addr <=  "0011000010010";
		Trees_din <= x"08ffd004";
		wait for Clk_period;
		Addr <=  "0011000010011";
		Trees_din <= x"00451869";
		wait for Clk_period;
		Addr <=  "0011000010100";
		Trees_din <= x"ff421869";
		wait for Clk_period;
		Addr <=  "0011000010101";
		Trees_din <= x"10007604";
		wait for Clk_period;
		Addr <=  "0011000010110";
		Trees_din <= x"ff2b1869";
		wait for Clk_period;
		Addr <=  "0011000010111";
		Trees_din <= x"e0ff4e04";
		wait for Clk_period;
		Addr <=  "0011000011000";
		Trees_din <= x"ffa01869";
		wait for Clk_period;
		Addr <=  "0011000011001";
		Trees_din <= x"00431869";
		wait for Clk_period;
		Addr <=  "0011000011010";
		Trees_din <= x"4400ba70";
		wait for Clk_period;
		Addr <=  "0011000011011";
		Trees_din <= x"d7008330";
		wait for Clk_period;
		Addr <=  "0011000011100";
		Trees_din <= x"fafea010";
		wait for Clk_period;
		Addr <=  "0011000011101";
		Trees_din <= x"f0ffb40c";
		wait for Clk_period;
		Addr <=  "0011000011110";
		Trees_din <= x"5a014e08";
		wait for Clk_period;
		Addr <=  "0011000011111";
		Trees_din <= x"db008204";
		wait for Clk_period;
		Addr <=  "0011000100000";
		Trees_din <= x"ff341975";
		wait for Clk_period;
		Addr <=  "0011000100001";
		Trees_din <= x"001e1975";
		wait for Clk_period;
		Addr <=  "0011000100010";
		Trees_din <= x"00511975";
		wait for Clk_period;
		Addr <=  "0011000100011";
		Trees_din <= x"00861975";
		wait for Clk_period;
		Addr <=  "0011000100100";
		Trees_din <= x"53ff7f10";
		wait for Clk_period;
		Addr <=  "0011000100101";
		Trees_din <= x"2bff3e08";
		wait for Clk_period;
		Addr <=  "0011000100110";
		Trees_din <= x"baffd304";
		wait for Clk_period;
		Addr <=  "0011000100111";
		Trees_din <= x"ffb11975";
		wait for Clk_period;
		Addr <=  "0011000101000";
		Trees_din <= x"002c1975";
		wait for Clk_period;
		Addr <=  "0011000101001";
		Trees_din <= x"99fe2404";
		wait for Clk_period;
		Addr <=  "0011000101010";
		Trees_din <= x"ffd51975";
		wait for Clk_period;
		Addr <=  "0011000101011";
		Trees_din <= x"00411975";
		wait for Clk_period;
		Addr <=  "0011000101100";
		Trees_din <= x"7eff0b08";
		wait for Clk_period;
		Addr <=  "0011000101101";
		Trees_din <= x"4bfe5204";
		wait for Clk_period;
		Addr <=  "0011000101110";
		Trees_din <= x"00601975";
		wait for Clk_period;
		Addr <=  "0011000101111";
		Trees_din <= x"fff01975";
		wait for Clk_period;
		Addr <=  "0011000110000";
		Trees_din <= x"b8ff1204";
		wait for Clk_period;
		Addr <=  "0011000110001";
		Trees_din <= x"ffb21975";
		wait for Clk_period;
		Addr <=  "0011000110010";
		Trees_din <= x"00431975";
		wait for Clk_period;
		Addr <=  "0011000110011";
		Trees_din <= x"21ff6820";
		wait for Clk_period;
		Addr <=  "0011000110100";
		Trees_din <= x"1fffbd10";
		wait for Clk_period;
		Addr <=  "0011000110101";
		Trees_din <= x"76ffbb08";
		wait for Clk_period;
		Addr <=  "0011000110110";
		Trees_din <= x"effee204";
		wait for Clk_period;
		Addr <=  "0011000110111";
		Trees_din <= x"ff721975";
		wait for Clk_period;
		Addr <=  "0011000111000";
		Trees_din <= x"00711975";
		wait for Clk_period;
		Addr <=  "0011000111001";
		Trees_din <= x"1afefd04";
		wait for Clk_period;
		Addr <=  "0011000111010";
		Trees_din <= x"ff761975";
		wait for Clk_period;
		Addr <=  "0011000111011";
		Trees_din <= x"00351975";
		wait for Clk_period;
		Addr <=  "0011000111100";
		Trees_din <= x"37ffec08";
		wait for Clk_period;
		Addr <=  "0011000111101";
		Trees_din <= x"16fe4a04";
		wait for Clk_period;
		Addr <=  "0011000111110";
		Trees_din <= x"ffed1975";
		wait for Clk_period;
		Addr <=  "0011000111111";
		Trees_din <= x"ff731975";
		wait for Clk_period;
		Addr <=  "0011001000000";
		Trees_din <= x"12ff8f04";
		wait for Clk_period;
		Addr <=  "0011001000001";
		Trees_din <= x"00931975";
		wait for Clk_period;
		Addr <=  "0011001000010";
		Trees_din <= x"ffb71975";
		wait for Clk_period;
		Addr <=  "0011001000011";
		Trees_din <= x"8fff2a10";
		wait for Clk_period;
		Addr <=  "0011001000100";
		Trees_din <= x"e9fe4a08";
		wait for Clk_period;
		Addr <=  "0011001000101";
		Trees_din <= x"cb001104";
		wait for Clk_period;
		Addr <=  "0011001000110";
		Trees_din <= x"ff7f1975";
		wait for Clk_period;
		Addr <=  "0011001000111";
		Trees_din <= x"00721975";
		wait for Clk_period;
		Addr <=  "0011001001000";
		Trees_din <= x"0400d204";
		wait for Clk_period;
		Addr <=  "0011001001001";
		Trees_din <= x"00351975";
		wait for Clk_period;
		Addr <=  "0011001001010";
		Trees_din <= x"ff8d1975";
		wait for Clk_period;
		Addr <=  "0011001001011";
		Trees_din <= x"ba002a08";
		wait for Clk_period;
		Addr <=  "0011001001100";
		Trees_din <= x"84ff6d04";
		wait for Clk_period;
		Addr <=  "0011001001101";
		Trees_din <= x"00191975";
		wait for Clk_period;
		Addr <=  "0011001001110";
		Trees_din <= x"ffb21975";
		wait for Clk_period;
		Addr <=  "0011001001111";
		Trees_din <= x"9aff5d04";
		wait for Clk_period;
		Addr <=  "0011001010000";
		Trees_din <= x"ff971975";
		wait for Clk_period;
		Addr <=  "0011001010001";
		Trees_din <= x"00911975";
		wait for Clk_period;
		Addr <=  "0011001010010";
		Trees_din <= x"dbffc410";
		wait for Clk_period;
		Addr <=  "0011001010011";
		Trees_din <= x"dfffc508";
		wait for Clk_period;
		Addr <=  "0011001010100";
		Trees_din <= x"05001204";
		wait for Clk_period;
		Addr <=  "0011001010101";
		Trees_din <= x"00331975";
		wait for Clk_period;
		Addr <=  "0011001010110";
		Trees_din <= x"ff711975";
		wait for Clk_period;
		Addr <=  "0011001010111";
		Trees_din <= x"6bfef304";
		wait for Clk_period;
		Addr <=  "0011001011000";
		Trees_din <= x"00931975";
		wait for Clk_period;
		Addr <=  "0011001011001";
		Trees_din <= x"00251975";
		wait for Clk_period;
		Addr <=  "0011001011010";
		Trees_din <= x"bbfed604";
		wait for Clk_period;
		Addr <=  "0011001011011";
		Trees_din <= x"00101975";
		wait for Clk_period;
		Addr <=  "0011001011100";
		Trees_din <= x"ff431975";
		wait for Clk_period;
		Addr <=  "0011001011101";
		Trees_din <= x"3fffb43c";
		wait for Clk_period;
		Addr <=  "0011001011110";
		Trees_din <= x"49ff620c";
		wait for Clk_period;
		Addr <=  "0011001011111";
		Trees_din <= x"26fff504";
		wait for Clk_period;
		Addr <=  "0011001100000";
		Trees_din <= x"005a1ab1";
		wait for Clk_period;
		Addr <=  "0011001100001";
		Trees_din <= x"06ff3b04";
		wait for Clk_period;
		Addr <=  "0011001100010";
		Trees_din <= x"ffd31ab1";
		wait for Clk_period;
		Addr <=  "0011001100011";
		Trees_din <= x"ff491ab1";
		wait for Clk_period;
		Addr <=  "0011001100100";
		Trees_din <= x"06fff520";
		wait for Clk_period;
		Addr <=  "0011001100101";
		Trees_din <= x"09001310";
		wait for Clk_period;
		Addr <=  "0011001100110";
		Trees_din <= x"33fef908";
		wait for Clk_period;
		Addr <=  "0011001100111";
		Trees_din <= x"cafe1004";
		wait for Clk_period;
		Addr <=  "0011001101000";
		Trees_din <= x"00571ab1";
		wait for Clk_period;
		Addr <=  "0011001101001";
		Trees_din <= x"ff821ab1";
		wait for Clk_period;
		Addr <=  "0011001101010";
		Trees_din <= x"c3ffcf04";
		wait for Clk_period;
		Addr <=  "0011001101011";
		Trees_din <= x"00161ab1";
		wait for Clk_period;
		Addr <=  "0011001101100";
		Trees_din <= x"00801ab1";
		wait for Clk_period;
		Addr <=  "0011001101101";
		Trees_din <= x"b0ff7508";
		wait for Clk_period;
		Addr <=  "0011001101110";
		Trees_din <= x"1bfffb04";
		wait for Clk_period;
		Addr <=  "0011001101111";
		Trees_din <= x"00671ab1";
		wait for Clk_period;
		Addr <=  "0011001110000";
		Trees_din <= x"ff831ab1";
		wait for Clk_period;
		Addr <=  "0011001110001";
		Trees_din <= x"99ff1904";
		wait for Clk_period;
		Addr <=  "0011001110010";
		Trees_din <= x"ffd11ab1";
		wait for Clk_period;
		Addr <=  "0011001110011";
		Trees_din <= x"ff281ab1";
		wait for Clk_period;
		Addr <=  "0011001110100";
		Trees_din <= x"9dffe408";
		wait for Clk_period;
		Addr <=  "0011001110101";
		Trees_din <= x"7bfed204";
		wait for Clk_period;
		Addr <=  "0011001110110";
		Trees_din <= x"ffe61ab1";
		wait for Clk_period;
		Addr <=  "0011001110111";
		Trees_din <= x"00b21ab1";
		wait for Clk_period;
		Addr <=  "0011001111000";
		Trees_din <= x"1dff1404";
		wait for Clk_period;
		Addr <=  "0011001111001";
		Trees_din <= x"00751ab1";
		wait for Clk_period;
		Addr <=  "0011001111010";
		Trees_din <= x"ff731ab1";
		wait for Clk_period;
		Addr <=  "0011001111011";
		Trees_din <= x"43ffa738";
		wait for Clk_period;
		Addr <=  "0011001111100";
		Trees_din <= x"24ff0d18";
		wait for Clk_period;
		Addr <=  "0011001111101";
		Trees_din <= x"56ff5108";
		wait for Clk_period;
		Addr <=  "0011001111110";
		Trees_din <= x"d6ffad04";
		wait for Clk_period;
		Addr <=  "0011001111111";
		Trees_din <= x"000a1ab1";
		wait for Clk_period;
		Addr <=  "0011010000000";
		Trees_din <= x"ff471ab1";
		wait for Clk_period;
		Addr <=  "0011010000001";
		Trees_din <= x"83ff5c08";
		wait for Clk_period;
		Addr <=  "0011010000010";
		Trees_din <= x"62fee304";
		wait for Clk_period;
		Addr <=  "0011010000011";
		Trees_din <= x"ff6f1ab1";
		wait for Clk_period;
		Addr <=  "0011010000100";
		Trees_din <= x"00401ab1";
		wait for Clk_period;
		Addr <=  "0011010000101";
		Trees_din <= x"eafed204";
		wait for Clk_period;
		Addr <=  "0011010000110";
		Trees_din <= x"00431ab1";
		wait for Clk_period;
		Addr <=  "0011010000111";
		Trees_din <= x"ff481ab1";
		wait for Clk_period;
		Addr <=  "0011010001000";
		Trees_din <= x"4cfeb310";
		wait for Clk_period;
		Addr <=  "0011010001001";
		Trees_din <= x"d700bf08";
		wait for Clk_period;
		Addr <=  "0011010001010";
		Trees_din <= x"24ff8104";
		wait for Clk_period;
		Addr <=  "0011010001011";
		Trees_din <= x"fff51ab1";
		wait for Clk_period;
		Addr <=  "0011010001100";
		Trees_din <= x"00501ab1";
		wait for Clk_period;
		Addr <=  "0011010001101";
		Trees_din <= x"ab007e04";
		wait for Clk_period;
		Addr <=  "0011010001110";
		Trees_din <= x"ff901ab1";
		wait for Clk_period;
		Addr <=  "0011010001111";
		Trees_din <= x"00741ab1";
		wait for Clk_period;
		Addr <=  "0011010010000";
		Trees_din <= x"bcff1808";
		wait for Clk_period;
		Addr <=  "0011010010001";
		Trees_din <= x"03ffb904";
		wait for Clk_period;
		Addr <=  "0011010010010";
		Trees_din <= x"fff91ab1";
		wait for Clk_period;
		Addr <=  "0011010010011";
		Trees_din <= x"ffb81ab1";
		wait for Clk_period;
		Addr <=  "0011010010100";
		Trees_din <= x"6d002904";
		wait for Clk_period;
		Addr <=  "0011010010101";
		Trees_din <= x"001f1ab1";
		wait for Clk_period;
		Addr <=  "0011010010110";
		Trees_din <= x"ffe91ab1";
		wait for Clk_period;
		Addr <=  "0011010010111";
		Trees_din <= x"06fed70c";
		wait for Clk_period;
		Addr <=  "0011010011000";
		Trees_din <= x"37ffce08";
		wait for Clk_period;
		Addr <=  "0011010011001";
		Trees_din <= x"cfffab04";
		wait for Clk_period;
		Addr <=  "0011010011010";
		Trees_din <= x"ffdd1ab1";
		wait for Clk_period;
		Addr <=  "0011010011011";
		Trees_din <= x"ff4a1ab1";
		wait for Clk_period;
		Addr <=  "0011010011100";
		Trees_din <= x"00361ab1";
		wait for Clk_period;
		Addr <=  "0011010011101";
		Trees_din <= x"0a00bc10";
		wait for Clk_period;
		Addr <=  "0011010011110";
		Trees_din <= x"ed005408";
		wait for Clk_period;
		Addr <=  "0011010011111";
		Trees_din <= x"f8ffe704";
		wait for Clk_period;
		Addr <=  "0011010100000";
		Trees_din <= x"fff11ab1";
		wait for Clk_period;
		Addr <=  "0011010100001";
		Trees_din <= x"00431ab1";
		wait for Clk_period;
		Addr <=  "0011010100010";
		Trees_din <= x"d2fed404";
		wait for Clk_period;
		Addr <=  "0011010100011";
		Trees_din <= x"00291ab1";
		wait for Clk_period;
		Addr <=  "0011010100100";
		Trees_din <= x"ff2c1ab1";
		wait for Clk_period;
		Addr <=  "0011010100101";
		Trees_din <= x"57ff2b08";
		wait for Clk_period;
		Addr <=  "0011010100110";
		Trees_din <= x"b7000904";
		wait for Clk_period;
		Addr <=  "0011010100111";
		Trees_din <= x"ff561ab1";
		wait for Clk_period;
		Addr <=  "0011010101000";
		Trees_din <= x"00291ab1";
		wait for Clk_period;
		Addr <=  "0011010101001";
		Trees_din <= x"65fef004";
		wait for Clk_period;
		Addr <=  "0011010101010";
		Trees_din <= x"ff921ab1";
		wait for Clk_period;
		Addr <=  "0011010101011";
		Trees_din <= x"00601ab1";
		wait for Clk_period;
		Addr <=  "0011010101100";
		Trees_din <= x"d5009d7c";
		wait for Clk_period;
		Addr <=  "0011010101101";
		Trees_din <= x"c8fff440";
		wait for Clk_period;
		Addr <=  "0011010101110";
		Trees_din <= x"50ff8420";
		wait for Clk_period;
		Addr <=  "0011010101111";
		Trees_din <= x"cf000710";
		wait for Clk_period;
		Addr <=  "0011010110000";
		Trees_din <= x"8eff6f08";
		wait for Clk_period;
		Addr <=  "0011010110001";
		Trees_din <= x"15ff0804";
		wait for Clk_period;
		Addr <=  "0011010110010";
		Trees_din <= x"006c1be5";
		wait for Clk_period;
		Addr <=  "0011010110011";
		Trees_din <= x"ff7d1be5";
		wait for Clk_period;
		Addr <=  "0011010110100";
		Trees_din <= x"81ff9804";
		wait for Clk_period;
		Addr <=  "0011010110101";
		Trees_din <= x"00151be5";
		wait for Clk_period;
		Addr <=  "0011010110110";
		Trees_din <= x"00611be5";
		wait for Clk_period;
		Addr <=  "0011010110111";
		Trees_din <= x"59ffdf08";
		wait for Clk_period;
		Addr <=  "0011010111000";
		Trees_din <= x"00ff5904";
		wait for Clk_period;
		Addr <=  "0011010111001";
		Trees_din <= x"fffb1be5";
		wait for Clk_period;
		Addr <=  "0011010111010";
		Trees_din <= x"ffa91be5";
		wait for Clk_period;
		Addr <=  "0011010111011";
		Trees_din <= x"89ffc904";
		wait for Clk_period;
		Addr <=  "0011010111100";
		Trees_din <= x"ffde1be5";
		wait for Clk_period;
		Addr <=  "0011010111101";
		Trees_din <= x"005b1be5";
		wait for Clk_period;
		Addr <=  "0011010111110";
		Trees_din <= x"93ff6d10";
		wait for Clk_period;
		Addr <=  "0011010111111";
		Trees_din <= x"49ffa608";
		wait for Clk_period;
		Addr <=  "0011011000000";
		Trees_din <= x"6d003c04";
		wait for Clk_period;
		Addr <=  "0011011000001";
		Trees_din <= x"00391be5";
		wait for Clk_period;
		Addr <=  "0011011000010";
		Trees_din <= x"ff781be5";
		wait for Clk_period;
		Addr <=  "0011011000011";
		Trees_din <= x"f8fff104";
		wait for Clk_period;
		Addr <=  "0011011000100";
		Trees_din <= x"00031be5";
		wait for Clk_period;
		Addr <=  "0011011000101";
		Trees_din <= x"00791be5";
		wait for Clk_period;
		Addr <=  "0011011000110";
		Trees_din <= x"44003008";
		wait for Clk_period;
		Addr <=  "0011011000111";
		Trees_din <= x"6affd304";
		wait for Clk_period;
		Addr <=  "0011011001000";
		Trees_din <= x"00431be5";
		wait for Clk_period;
		Addr <=  "0011011001001";
		Trees_din <= x"ffd41be5";
		wait for Clk_period;
		Addr <=  "0011011001010";
		Trees_din <= x"f6fea704";
		wait for Clk_period;
		Addr <=  "0011011001011";
		Trees_din <= x"003e1be5";
		wait for Clk_period;
		Addr <=  "0011011001100";
		Trees_din <= x"ffa21be5";
		wait for Clk_period;
		Addr <=  "0011011001101";
		Trees_din <= x"27003c20";
		wait for Clk_period;
		Addr <=  "0011011001110";
		Trees_din <= x"65ffeb10";
		wait for Clk_period;
		Addr <=  "0011011001111";
		Trees_din <= x"0dffe308";
		wait for Clk_period;
		Addr <=  "0011011010000";
		Trees_din <= x"b2ffd704";
		wait for Clk_period;
		Addr <=  "0011011010001";
		Trees_din <= x"ffcc1be5";
		wait for Clk_period;
		Addr <=  "0011011010010";
		Trees_din <= x"00031be5";
		wait for Clk_period;
		Addr <=  "0011011010011";
		Trees_din <= x"76ff6904";
		wait for Clk_period;
		Addr <=  "0011011010100";
		Trees_din <= x"ffc31be5";
		wait for Clk_period;
		Addr <=  "0011011010101";
		Trees_din <= x"00381be5";
		wait for Clk_period;
		Addr <=  "0011011010110";
		Trees_din <= x"7dffe208";
		wait for Clk_period;
		Addr <=  "0011011010111";
		Trees_din <= x"e3fe5e04";
		wait for Clk_period;
		Addr <=  "0011011011000";
		Trees_din <= x"00051be5";
		wait for Clk_period;
		Addr <=  "0011011011001";
		Trees_din <= x"00a41be5";
		wait for Clk_period;
		Addr <=  "0011011011010";
		Trees_din <= x"f8009c04";
		wait for Clk_period;
		Addr <=  "0011011011011";
		Trees_din <= x"00431be5";
		wait for Clk_period;
		Addr <=  "0011011011100";
		Trees_din <= x"ff921be5";
		wait for Clk_period;
		Addr <=  "0011011011101";
		Trees_din <= x"5a00f510";
		wait for Clk_period;
		Addr <=  "0011011011110";
		Trees_din <= x"5bffa108";
		wait for Clk_period;
		Addr <=  "0011011011111";
		Trees_din <= x"59002e04";
		wait for Clk_period;
		Addr <=  "0011011100000";
		Trees_din <= x"ff801be5";
		wait for Clk_period;
		Addr <=  "0011011100001";
		Trees_din <= x"00081be5";
		wait for Clk_period;
		Addr <=  "0011011100010";
		Trees_din <= x"5dffeb04";
		wait for Clk_period;
		Addr <=  "0011011100011";
		Trees_din <= x"ffd61be5";
		wait for Clk_period;
		Addr <=  "0011011100100";
		Trees_din <= x"008a1be5";
		wait for Clk_period;
		Addr <=  "0011011100101";
		Trees_din <= x"cafddb04";
		wait for Clk_period;
		Addr <=  "0011011100110";
		Trees_din <= x"ff831be5";
		wait for Clk_period;
		Addr <=  "0011011100111";
		Trees_din <= x"93ff7f04";
		wait for Clk_period;
		Addr <=  "0011011101000";
		Trees_din <= x"00a11be5";
		wait for Clk_period;
		Addr <=  "0011011101001";
		Trees_din <= x"ffd91be5";
		wait for Clk_period;
		Addr <=  "0011011101010";
		Trees_din <= x"78fee00c";
		wait for Clk_period;
		Addr <=  "0011011101011";
		Trees_din <= x"fdff5c08";
		wait for Clk_period;
		Addr <=  "0011011101100";
		Trees_din <= x"b4ff3004";
		wait for Clk_period;
		Addr <=  "0011011101101";
		Trees_din <= x"00231be5";
		wait for Clk_period;
		Addr <=  "0011011101110";
		Trees_din <= x"00931be5";
		wait for Clk_period;
		Addr <=  "0011011101111";
		Trees_din <= x"ffc21be5";
		wait for Clk_period;
		Addr <=  "0011011110000";
		Trees_din <= x"1dfe8f08";
		wait for Clk_period;
		Addr <=  "0011011110001";
		Trees_din <= x"f7ff0304";
		wait for Clk_period;
		Addr <=  "0011011110010";
		Trees_din <= x"00611be5";
		wait for Clk_period;
		Addr <=  "0011011110011";
		Trees_din <= x"ffed1be5";
		wait for Clk_period;
		Addr <=  "0011011110100";
		Trees_din <= x"04003704";
		wait for Clk_period;
		Addr <=  "0011011110101";
		Trees_din <= x"002b1be5";
		wait for Clk_period;
		Addr <=  "0011011110110";
		Trees_din <= x"8fff9504";
		wait for Clk_period;
		Addr <=  "0011011110111";
		Trees_din <= x"ff4e1be5";
		wait for Clk_period;
		Addr <=  "0011011111000";
		Trees_din <= x"ffc71be5";
		wait for Clk_period;
		Addr <=  "0011011111001";
		Trees_din <= x"40005868";
		wait for Clk_period;
		Addr <=  "0011011111010";
		Trees_din <= x"cafdaa28";
		wait for Clk_period;
		Addr <=  "0011011111011";
		Trees_din <= x"7dffef14";
		wait for Clk_period;
		Addr <=  "0011011111100";
		Trees_din <= x"5bffdb10";
		wait for Clk_period;
		Addr <=  "0011011111101";
		Trees_din <= x"03ff5d08";
		wait for Clk_period;
		Addr <=  "0011011111110";
		Trees_din <= x"b3ff0504";
		wait for Clk_period;
		Addr <=  "0011011111111";
		Trees_din <= x"ffd81d59";
		wait for Clk_period;
		Addr <=  "0011100000000";
		Trees_din <= x"008c1d59";
		wait for Clk_period;
		Addr <=  "0011100000001";
		Trees_din <= x"32feef04";
		wait for Clk_period;
		Addr <=  "0011100000010";
		Trees_din <= x"fff71d59";
		wait for Clk_period;
		Addr <=  "0011100000011";
		Trees_din <= x"ff5f1d59";
		wait for Clk_period;
		Addr <=  "0011100000100";
		Trees_din <= x"00b51d59";
		wait for Clk_period;
		Addr <=  "0011100000101";
		Trees_din <= x"07ffc208";
		wait for Clk_period;
		Addr <=  "0011100000110";
		Trees_din <= x"10ffe504";
		wait for Clk_period;
		Addr <=  "0011100000111";
		Trees_din <= x"005c1d59";
		wait for Clk_period;
		Addr <=  "0011100001000";
		Trees_din <= x"ffb41d59";
		wait for Clk_period;
		Addr <=  "0011100001001";
		Trees_din <= x"71ffcb08";
		wait for Clk_period;
		Addr <=  "0011100001010";
		Trees_din <= x"ad000304";
		wait for Clk_period;
		Addr <=  "0011100001011";
		Trees_din <= x"ff381d59";
		wait for Clk_period;
		Addr <=  "0011100001100";
		Trees_din <= x"00161d59";
		wait for Clk_period;
		Addr <=  "0011100001101";
		Trees_din <= x"003b1d59";
		wait for Clk_period;
		Addr <=  "0011100001110";
		Trees_din <= x"d7007c20";
		wait for Clk_period;
		Addr <=  "0011100001111";
		Trees_din <= x"fafea010";
		wait for Clk_period;
		Addr <=  "0011100010000";
		Trees_din <= x"f201a808";
		wait for Clk_period;
		Addr <=  "0011100010001";
		Trees_din <= x"00ff4804";
		wait for Clk_period;
		Addr <=  "0011100010010";
		Trees_din <= x"00591d59";
		wait for Clk_period;
		Addr <=  "0011100010011";
		Trees_din <= x"fffc1d59";
		wait for Clk_period;
		Addr <=  "0011100010100";
		Trees_din <= x"e4fe7504";
		wait for Clk_period;
		Addr <=  "0011100010101";
		Trees_din <= x"000e1d59";
		wait for Clk_period;
		Addr <=  "0011100010110";
		Trees_din <= x"ff431d59";
		wait for Clk_period;
		Addr <=  "0011100010111";
		Trees_din <= x"63ff9f08";
		wait for Clk_period;
		Addr <=  "0011100011000";
		Trees_din <= x"bcfeff04";
		wait for Clk_period;
		Addr <=  "0011100011001";
		Trees_din <= x"000f1d59";
		wait for Clk_period;
		Addr <=  "0011100011010";
		Trees_din <= x"00451d59";
		wait for Clk_period;
		Addr <=  "0011100011011";
		Trees_din <= x"f8009904";
		wait for Clk_period;
		Addr <=  "0011100011100";
		Trees_din <= x"00181d59";
		wait for Clk_period;
		Addr <=  "0011100011101";
		Trees_din <= x"ffca1d59";
		wait for Clk_period;
		Addr <=  "0011100011110";
		Trees_din <= x"21ffd310";
		wait for Clk_period;
		Addr <=  "0011100011111";
		Trees_din <= x"a0fe3d08";
		wait for Clk_period;
		Addr <=  "0011100100000";
		Trees_din <= x"0efe4004";
		wait for Clk_period;
		Addr <=  "0011100100001";
		Trees_din <= x"ffcd1d59";
		wait for Clk_period;
		Addr <=  "0011100100010";
		Trees_din <= x"005f1d59";
		wait for Clk_period;
		Addr <=  "0011100100011";
		Trees_din <= x"3fff9404";
		wait for Clk_period;
		Addr <=  "0011100100100";
		Trees_din <= x"005e1d59";
		wait for Clk_period;
		Addr <=  "0011100100101";
		Trees_din <= x"ffcc1d59";
		wait for Clk_period;
		Addr <=  "0011100100110";
		Trees_din <= x"1eff7108";
		wait for Clk_period;
		Addr <=  "0011100100111";
		Trees_din <= x"06ff9e04";
		wait for Clk_period;
		Addr <=  "0011100101000";
		Trees_din <= x"00251d59";
		wait for Clk_period;
		Addr <=  "0011100101001";
		Trees_din <= x"ff9f1d59";
		wait for Clk_period;
		Addr <=  "0011100101010";
		Trees_din <= x"ce009104";
		wait for Clk_period;
		Addr <=  "0011100101011";
		Trees_din <= x"00491d59";
		wait for Clk_period;
		Addr <=  "0011100101100";
		Trees_din <= x"ff3f1d59";
		wait for Clk_period;
		Addr <=  "0011100101101";
		Trees_din <= x"1aff142c";
		wait for Clk_period;
		Addr <=  "0011100101110";
		Trees_din <= x"aeff8d18";
		wait for Clk_period;
		Addr <=  "0011100101111";
		Trees_din <= x"34ff7d08";
		wait for Clk_period;
		Addr <=  "0011100110000";
		Trees_din <= x"11ff7c04";
		wait for Clk_period;
		Addr <=  "0011100110001";
		Trees_din <= x"00971d59";
		wait for Clk_period;
		Addr <=  "0011100110010";
		Trees_din <= x"ffda1d59";
		wait for Clk_period;
		Addr <=  "0011100110011";
		Trees_din <= x"0bff2508";
		wait for Clk_period;
		Addr <=  "0011100110100";
		Trees_din <= x"a9ffa604";
		wait for Clk_period;
		Addr <=  "0011100110101";
		Trees_din <= x"008d1d59";
		wait for Clk_period;
		Addr <=  "0011100110110";
		Trees_din <= x"ffa71d59";
		wait for Clk_period;
		Addr <=  "0011100110111";
		Trees_din <= x"4bfe1004";
		wait for Clk_period;
		Addr <=  "0011100111000";
		Trees_din <= x"00621d59";
		wait for Clk_period;
		Addr <=  "0011100111001";
		Trees_din <= x"ff861d59";
		wait for Clk_period;
		Addr <=  "0011100111010";
		Trees_din <= x"51002a0c";
		wait for Clk_period;
		Addr <=  "0011100111011";
		Trees_din <= x"52ff0404";
		wait for Clk_period;
		Addr <=  "0011100111100";
		Trees_din <= x"ffca1d59";
		wait for Clk_period;
		Addr <=  "0011100111101";
		Trees_din <= x"18ff5204";
		wait for Clk_period;
		Addr <=  "0011100111110";
		Trees_din <= x"00191d59";
		wait for Clk_period;
		Addr <=  "0011100111111";
		Trees_din <= x"00a01d59";
		wait for Clk_period;
		Addr <=  "0011101000000";
		Trees_din <= x"c8003804";
		wait for Clk_period;
		Addr <=  "0011101000001";
		Trees_din <= x"ff891d59";
		wait for Clk_period;
		Addr <=  "0011101000010";
		Trees_din <= x"000c1d59";
		wait for Clk_period;
		Addr <=  "0011101000011";
		Trees_din <= x"11ffab1c";
		wait for Clk_period;
		Addr <=  "0011101000100";
		Trees_din <= x"8effa90c";
		wait for Clk_period;
		Addr <=  "0011101000101";
		Trees_din <= x"28ff6508";
		wait for Clk_period;
		Addr <=  "0011101000110";
		Trees_din <= x"aafee204";
		wait for Clk_period;
		Addr <=  "0011101000111";
		Trees_din <= x"00281d59";
		wait for Clk_period;
		Addr <=  "0011101001000";
		Trees_din <= x"ff531d59";
		wait for Clk_period;
		Addr <=  "0011101001001";
		Trees_din <= x"00691d59";
		wait for Clk_period;
		Addr <=  "0011101001010";
		Trees_din <= x"48ff5308";
		wait for Clk_period;
		Addr <=  "0011101001011";
		Trees_din <= x"c0ff2504";
		wait for Clk_period;
		Addr <=  "0011101001100";
		Trees_din <= x"00221d59";
		wait for Clk_period;
		Addr <=  "0011101001101";
		Trees_din <= x"ff741d59";
		wait for Clk_period;
		Addr <=  "0011101001110";
		Trees_din <= x"87ff4b04";
		wait for Clk_period;
		Addr <=  "0011101001111";
		Trees_din <= x"ffff1d59";
		wait for Clk_period;
		Addr <=  "0011101010000";
		Trees_din <= x"00951d59";
		wait for Clk_period;
		Addr <=  "0011101010001";
		Trees_din <= x"53ff6b04";
		wait for Clk_period;
		Addr <=  "0011101010010";
		Trees_din <= x"00321d59";
		wait for Clk_period;
		Addr <=  "0011101010011";
		Trees_din <= x"e7ffd304";
		wait for Clk_period;
		Addr <=  "0011101010100";
		Trees_din <= x"ff501d59";
		wait for Clk_period;
		Addr <=  "0011101010101";
		Trees_din <= x"fff61d59";
		wait for Clk_period;
		Addr <=  "0011101010110";
		Trees_din <= x"49ffa558";
		wait for Clk_period;
		Addr <=  "0011101010111";
		Trees_din <= x"0bff5a24";
		wait for Clk_period;
		Addr <=  "0011101011000";
		Trees_din <= x"daff4d08";
		wait for Clk_period;
		Addr <=  "0011101011001";
		Trees_din <= x"faff6e04";
		wait for Clk_period;
		Addr <=  "0011101011010";
		Trees_din <= x"ff691ef5";
		wait for Clk_period;
		Addr <=  "0011101011011";
		Trees_din <= x"000e1ef5";
		wait for Clk_period;
		Addr <=  "0011101011100";
		Trees_din <= x"42ff9a0c";
		wait for Clk_period;
		Addr <=  "0011101011101";
		Trees_din <= x"e5fe5704";
		wait for Clk_period;
		Addr <=  "0011101011110";
		Trees_din <= x"ffbd1ef5";
		wait for Clk_period;
		Addr <=  "0011101011111";
		Trees_din <= x"2bfeec04";
		wait for Clk_period;
		Addr <=  "0011101100000";
		Trees_din <= x"00071ef5";
		wait for Clk_period;
		Addr <=  "0011101100001";
		Trees_din <= x"00a61ef5";
		wait for Clk_period;
		Addr <=  "0011101100010";
		Trees_din <= x"35ff0608";
		wait for Clk_period;
		Addr <=  "0011101100011";
		Trees_din <= x"56ffe804";
		wait for Clk_period;
		Addr <=  "0011101100100";
		Trees_din <= x"ff921ef5";
		wait for Clk_period;
		Addr <=  "0011101100101";
		Trees_din <= x"00691ef5";
		wait for Clk_period;
		Addr <=  "0011101100110";
		Trees_din <= x"d6007d04";
		wait for Clk_period;
		Addr <=  "0011101100111";
		Trees_din <= x"00931ef5";
		wait for Clk_period;
		Addr <=  "0011101101000";
		Trees_din <= x"00091ef5";
		wait for Clk_period;
		Addr <=  "0011101101001";
		Trees_din <= x"7eff2118";
		wait for Clk_period;
		Addr <=  "0011101101010";
		Trees_din <= x"59008d10";
		wait for Clk_period;
		Addr <=  "0011101101011";
		Trees_din <= x"e1ffba08";
		wait for Clk_period;
		Addr <=  "0011101101100";
		Trees_din <= x"d6009504";
		wait for Clk_period;
		Addr <=  "0011101101101";
		Trees_din <= x"ffc81ef5";
		wait for Clk_period;
		Addr <=  "0011101101110";
		Trees_din <= x"003f1ef5";
		wait for Clk_period;
		Addr <=  "0011101101111";
		Trees_din <= x"52ff6504";
		wait for Clk_period;
		Addr <=  "0011101110000";
		Trees_din <= x"ff831ef5";
		wait for Clk_period;
		Addr <=  "0011101110001";
		Trees_din <= x"ffe11ef5";
		wait for Clk_period;
		Addr <=  "0011101110010";
		Trees_din <= x"36ff8f04";
		wait for Clk_period;
		Addr <=  "0011101110011";
		Trees_din <= x"009f1ef5";
		wait for Clk_period;
		Addr <=  "0011101110100";
		Trees_din <= x"ffb81ef5";
		wait for Clk_period;
		Addr <=  "0011101110101";
		Trees_din <= x"0400a410";
		wait for Clk_period;
		Addr <=  "0011101110110";
		Trees_din <= x"12fff608";
		wait for Clk_period;
		Addr <=  "0011101110111";
		Trees_din <= x"93ffe104";
		wait for Clk_period;
		Addr <=  "0011101111000";
		Trees_din <= x"00561ef5";
		wait for Clk_period;
		Addr <=  "0011101111001";
		Trees_din <= x"ffab1ef5";
		wait for Clk_period;
		Addr <=  "0011101111010";
		Trees_din <= x"b8ff8d04";
		wait for Clk_period;
		Addr <=  "0011101111011";
		Trees_din <= x"ff621ef5";
		wait for Clk_period;
		Addr <=  "0011101111100";
		Trees_din <= x"00311ef5";
		wait for Clk_period;
		Addr <=  "0011101111101";
		Trees_din <= x"15ff4a04";
		wait for Clk_period;
		Addr <=  "0011101111110";
		Trees_din <= x"00681ef5";
		wait for Clk_period;
		Addr <=  "0011101111111";
		Trees_din <= x"79ff0104";
		wait for Clk_period;
		Addr <=  "0011110000000";
		Trees_din <= x"ffcc1ef5";
		wait for Clk_period;
		Addr <=  "0011110000001";
		Trees_din <= x"ff3f1ef5";
		wait for Clk_period;
		Addr <=  "0011110000010";
		Trees_din <= x"dc003c40";
		wait for Clk_period;
		Addr <=  "0011110000011";
		Trees_din <= x"da006520";
		wait for Clk_period;
		Addr <=  "0011110000100";
		Trees_din <= x"3eff8210";
		wait for Clk_period;
		Addr <=  "0011110000101";
		Trees_din <= x"4400b408";
		wait for Clk_period;
		Addr <=  "0011110000110";
		Trees_din <= x"0d002d04";
		wait for Clk_period;
		Addr <=  "0011110000111";
		Trees_din <= x"00241ef5";
		wait for Clk_period;
		Addr <=  "0011110001000";
		Trees_din <= x"006a1ef5";
		wait for Clk_period;
		Addr <=  "0011110001001";
		Trees_din <= x"c9ffb004";
		wait for Clk_period;
		Addr <=  "0011110001010";
		Trees_din <= x"002a1ef5";
		wait for Clk_period;
		Addr <=  "0011110001011";
		Trees_din <= x"ff571ef5";
		wait for Clk_period;
		Addr <=  "0011110001100";
		Trees_din <= x"9bff4b08";
		wait for Clk_period;
		Addr <=  "0011110001101";
		Trees_din <= x"afff0604";
		wait for Clk_period;
		Addr <=  "0011110001110";
		Trees_din <= x"00631ef5";
		wait for Clk_period;
		Addr <=  "0011110001111";
		Trees_din <= x"ffc81ef5";
		wait for Clk_period;
		Addr <=  "0011110010000";
		Trees_din <= x"6bfe5f04";
		wait for Clk_period;
		Addr <=  "0011110010001";
		Trees_din <= x"ff861ef5";
		wait for Clk_period;
		Addr <=  "0011110010010";
		Trees_din <= x"00211ef5";
		wait for Clk_period;
		Addr <=  "0011110010011";
		Trees_din <= x"6fff8f10";
		wait for Clk_period;
		Addr <=  "0011110010100";
		Trees_din <= x"0cfe7008";
		wait for Clk_period;
		Addr <=  "0011110010101";
		Trees_din <= x"1afefb04";
		wait for Clk_period;
		Addr <=  "0011110010110";
		Trees_din <= x"ff9c1ef5";
		wait for Clk_period;
		Addr <=  "0011110010111";
		Trees_din <= x"00651ef5";
		wait for Clk_period;
		Addr <=  "0011110011000";
		Trees_din <= x"6cfed104";
		wait for Clk_period;
		Addr <=  "0011110011001";
		Trees_din <= x"00251ef5";
		wait for Clk_period;
		Addr <=  "0011110011010";
		Trees_din <= x"ff501ef5";
		wait for Clk_period;
		Addr <=  "0011110011011";
		Trees_din <= x"9ffeea08";
		wait for Clk_period;
		Addr <=  "0011110011100";
		Trees_din <= x"d5fff904";
		wait for Clk_period;
		Addr <=  "0011110011101";
		Trees_din <= x"000f1ef5";
		wait for Clk_period;
		Addr <=  "0011110011110";
		Trees_din <= x"ff561ef5";
		wait for Clk_period;
		Addr <=  "0011110011111";
		Trees_din <= x"9bfecd04";
		wait for Clk_period;
		Addr <=  "0011110100000";
		Trees_din <= x"ff871ef5";
		wait for Clk_period;
		Addr <=  "0011110100001";
		Trees_din <= x"00351ef5";
		wait for Clk_period;
		Addr <=  "0011110100010";
		Trees_din <= x"1dfeb118";
		wait for Clk_period;
		Addr <=  "0011110100011";
		Trees_din <= x"b7ffa70c";
		wait for Clk_period;
		Addr <=  "0011110100100";
		Trees_din <= x"43ffb008";
		wait for Clk_period;
		Addr <=  "0011110100101";
		Trees_din <= x"65ff9a04";
		wait for Clk_period;
		Addr <=  "0011110100110";
		Trees_din <= x"ff5a1ef5";
		wait for Clk_period;
		Addr <=  "0011110100111";
		Trees_din <= x"003a1ef5";
		wait for Clk_period;
		Addr <=  "0011110101000";
		Trees_din <= x"00671ef5";
		wait for Clk_period;
		Addr <=  "0011110101001";
		Trees_din <= x"19ff0404";
		wait for Clk_period;
		Addr <=  "0011110101010";
		Trees_din <= x"ff811ef5";
		wait for Clk_period;
		Addr <=  "0011110101011";
		Trees_din <= x"0dfef904";
		wait for Clk_period;
		Addr <=  "0011110101100";
		Trees_din <= x"ffd41ef5";
		wait for Clk_period;
		Addr <=  "0011110101101";
		Trees_din <= x"009c1ef5";
		wait for Clk_period;
		Addr <=  "0011110101110";
		Trees_din <= x"60ff6c10";
		wait for Clk_period;
		Addr <=  "0011110101111";
		Trees_din <= x"72005508";
		wait for Clk_period;
		Addr <=  "0011110110000";
		Trees_din <= x"e1000004";
		wait for Clk_period;
		Addr <=  "0011110110001";
		Trees_din <= x"00471ef5";
		wait for Clk_period;
		Addr <=  "0011110110010";
		Trees_din <= x"ffbf1ef5";
		wait for Clk_period;
		Addr <=  "0011110110011";
		Trees_din <= x"b3fe7b04";
		wait for Clk_period;
		Addr <=  "0011110110100";
		Trees_din <= x"00441ef5";
		wait for Clk_period;
		Addr <=  "0011110110101";
		Trees_din <= x"ff691ef5";
		wait for Clk_period;
		Addr <=  "0011110110110";
		Trees_din <= x"c9ff9208";
		wait for Clk_period;
		Addr <=  "0011110110111";
		Trees_din <= x"ddff2104";
		wait for Clk_period;
		Addr <=  "0011110111000";
		Trees_din <= x"ff9a1ef5";
		wait for Clk_period;
		Addr <=  "0011110111001";
		Trees_din <= x"00511ef5";
		wait for Clk_period;
		Addr <=  "0011110111010";
		Trees_din <= x"1aff5a04";
		wait for Clk_period;
		Addr <=  "0011110111011";
		Trees_din <= x"ff6c1ef5";
		wait for Clk_period;
		Addr <=  "0011110111100";
		Trees_din <= x"00531ef5";
		wait for Clk_period;
		Addr <=  "0011110111101";
		Trees_din <= x"f5007e80";
		wait for Clk_period;
		Addr <=  "0011110111110";
		Trees_din <= x"afff5640";
		wait for Clk_period;
		Addr <=  "0011110111111";
		Trees_din <= x"2fff6420";
		wait for Clk_period;
		Addr <=  "0011111000000";
		Trees_din <= x"e5fe9110";
		wait for Clk_period;
		Addr <=  "0011111000001";
		Trees_din <= x"10ff5108";
		wait for Clk_period;
		Addr <=  "0011111000010";
		Trees_din <= x"82ff3404";
		wait for Clk_period;
		Addr <=  "0011111000011";
		Trees_din <= x"00652049";
		wait for Clk_period;
		Addr <=  "0011111000100";
		Trees_din <= x"ffde2049";
		wait for Clk_period;
		Addr <=  "0011111000101";
		Trees_din <= x"35fff904";
		wait for Clk_period;
		Addr <=  "0011111000110";
		Trees_din <= x"ff972049";
		wait for Clk_period;
		Addr <=  "0011111000111";
		Trees_din <= x"00602049";
		wait for Clk_period;
		Addr <=  "0011111001000";
		Trees_din <= x"3cff3e08";
		wait for Clk_period;
		Addr <=  "0011111001001";
		Trees_din <= x"64fef704";
		wait for Clk_period;
		Addr <=  "0011111001010";
		Trees_din <= x"00602049";
		wait for Clk_period;
		Addr <=  "0011111001011";
		Trees_din <= x"ffdc2049";
		wait for Clk_period;
		Addr <=  "0011111001100";
		Trees_din <= x"3ffffc04";
		wait for Clk_period;
		Addr <=  "0011111001101";
		Trees_din <= x"00ae2049";
		wait for Clk_period;
		Addr <=  "0011111001110";
		Trees_din <= x"002a2049";
		wait for Clk_period;
		Addr <=  "0011111001111";
		Trees_din <= x"58ff9710";
		wait for Clk_period;
		Addr <=  "0011111010000";
		Trees_din <= x"96ff9308";
		wait for Clk_period;
		Addr <=  "0011111010001";
		Trees_din <= x"2fffa704";
		wait for Clk_period;
		Addr <=  "0011111010010";
		Trees_din <= x"ff692049";
		wait for Clk_period;
		Addr <=  "0011111010011";
		Trees_din <= x"ffcd2049";
		wait for Clk_period;
		Addr <=  "0011111010100";
		Trees_din <= x"b3ff0704";
		wait for Clk_period;
		Addr <=  "0011111010101";
		Trees_din <= x"ffa12049";
		wait for Clk_period;
		Addr <=  "0011111010110";
		Trees_din <= x"00572049";
		wait for Clk_period;
		Addr <=  "0011111010111";
		Trees_din <= x"8bfff808";
		wait for Clk_period;
		Addr <=  "0011111011000";
		Trees_din <= x"16ff6604";
		wait for Clk_period;
		Addr <=  "0011111011001";
		Trees_din <= x"ff7b2049";
		wait for Clk_period;
		Addr <=  "0011111011010";
		Trees_din <= x"00242049";
		wait for Clk_period;
		Addr <=  "0011111011011";
		Trees_din <= x"8c000e04";
		wait for Clk_period;
		Addr <=  "0011111011100";
		Trees_din <= x"009d2049";
		wait for Clk_period;
		Addr <=  "0011111011101";
		Trees_din <= x"ffe62049";
		wait for Clk_period;
		Addr <=  "0011111011110";
		Trees_din <= x"ddfede20";
		wait for Clk_period;
		Addr <=  "0011111011111";
		Trees_din <= x"64ff0b10";
		wait for Clk_period;
		Addr <=  "0011111100000";
		Trees_din <= x"e6ff5308";
		wait for Clk_period;
		Addr <=  "0011111100001";
		Trees_din <= x"2a00e804";
		wait for Clk_period;
		Addr <=  "0011111100010";
		Trees_din <= x"007b2049";
		wait for Clk_period;
		Addr <=  "0011111100011";
		Trees_din <= x"ff9c2049";
		wait for Clk_period;
		Addr <=  "0011111100100";
		Trees_din <= x"59007d04";
		wait for Clk_period;
		Addr <=  "0011111100101";
		Trees_din <= x"ff9e2049";
		wait for Clk_period;
		Addr <=  "0011111100110";
		Trees_din <= x"006e2049";
		wait for Clk_period;
		Addr <=  "0011111100111";
		Trees_din <= x"c9ff5708";
		wait for Clk_period;
		Addr <=  "0011111101000";
		Trees_din <= x"40004104";
		wait for Clk_period;
		Addr <=  "0011111101001";
		Trees_din <= x"00992049";
		wait for Clk_period;
		Addr <=  "0011111101010";
		Trees_din <= x"ffe12049";
		wait for Clk_period;
		Addr <=  "0011111101011";
		Trees_din <= x"64ffc404";
		wait for Clk_period;
		Addr <=  "0011111101100";
		Trees_din <= x"00072049";
		wait for Clk_period;
		Addr <=  "0011111101101";
		Trees_din <= x"ff9c2049";
		wait for Clk_period;
		Addr <=  "0011111101110";
		Trees_din <= x"71001310";
		wait for Clk_period;
		Addr <=  "0011111101111";
		Trees_din <= x"e9fe2708";
		wait for Clk_period;
		Addr <=  "0011111110000";
		Trees_din <= x"8dfe5404";
		wait for Clk_period;
		Addr <=  "0011111110001";
		Trees_din <= x"000f2049";
		wait for Clk_period;
		Addr <=  "0011111110010";
		Trees_din <= x"ff6e2049";
		wait for Clk_period;
		Addr <=  "0011111110011";
		Trees_din <= x"5a014904";
		wait for Clk_period;
		Addr <=  "0011111110100";
		Trees_din <= x"00142049";
		wait for Clk_period;
		Addr <=  "0011111110101";
		Trees_din <= x"00642049";
		wait for Clk_period;
		Addr <=  "0011111110110";
		Trees_din <= x"a8ffc308";
		wait for Clk_period;
		Addr <=  "0011111110111";
		Trees_din <= x"75ffde04";
		wait for Clk_period;
		Addr <=  "0011111111000";
		Trees_din <= x"fffa2049";
		wait for Clk_period;
		Addr <=  "0011111111001";
		Trees_din <= x"ff462049";
		wait for Clk_period;
		Addr <=  "0011111111010";
		Trees_din <= x"9bff2104";
		wait for Clk_period;
		Addr <=  "0011111111011";
		Trees_din <= x"ffb32049";
		wait for Clk_period;
		Addr <=  "0011111111100";
		Trees_din <= x"00802049";
		wait for Clk_period;
		Addr <=  "0011111111101";
		Trees_din <= x"2dff4320";
		wait for Clk_period;
		Addr <=  "0011111111110";
		Trees_din <= x"5400ec18";
		wait for Clk_period;
		Addr <=  "0011111111111";
		Trees_din <= x"2aff860c";
		wait for Clk_period;
		Addr <=  "0100000000000";
		Trees_din <= x"4dfe3104";
		wait for Clk_period;
		Addr <=  "0100000000001";
		Trees_din <= x"ff872049";
		wait for Clk_period;
		Addr <=  "0100000000010";
		Trees_din <= x"9affee04";
		wait for Clk_period;
		Addr <=  "0100000000011";
		Trees_din <= x"00712049";
		wait for Clk_period;
		Addr <=  "0100000000100";
		Trees_din <= x"00182049";
		wait for Clk_period;
		Addr <=  "0100000000101";
		Trees_din <= x"a5fe9104";
		wait for Clk_period;
		Addr <=  "0100000000110";
		Trees_din <= x"ffdc2049";
		wait for Clk_period;
		Addr <=  "0100000000111";
		Trees_din <= x"82ffcf04";
		wait for Clk_period;
		Addr <=  "0100000001000";
		Trees_din <= x"00a02049";
		wait for Clk_period;
		Addr <=  "0100000001001";
		Trees_din <= x"fff82049";
		wait for Clk_period;
		Addr <=  "0100000001010";
		Trees_din <= x"a5fed004";
		wait for Clk_period;
		Addr <=  "0100000001011";
		Trees_din <= x"00622049";
		wait for Clk_period;
		Addr <=  "0100000001100";
		Trees_din <= x"ff422049";
		wait for Clk_period;
		Addr <=  "0100000001101";
		Trees_din <= x"e3fe9d08";
		wait for Clk_period;
		Addr <=  "0100000001110";
		Trees_din <= x"34ffd404";
		wait for Clk_period;
		Addr <=  "0100000001111";
		Trees_din <= x"ffe12049";
		wait for Clk_period;
		Addr <=  "0100000010000";
		Trees_din <= x"ff792049";
		wait for Clk_period;
		Addr <=  "0100000010001";
		Trees_din <= x"00192049";
		wait for Clk_period;
		Addr <=  "0100000010010";
		Trees_din <= x"b6ff7274";
		wait for Clk_period;
		Addr <=  "0100000010011";
		Trees_din <= x"9bff3d40";
		wait for Clk_period;
		Addr <=  "0100000010100";
		Trees_din <= x"3f002220";
		wait for Clk_period;
		Addr <=  "0100000010101";
		Trees_din <= x"e0feb810";
		wait for Clk_period;
		Addr <=  "0100000010110";
		Trees_din <= x"76ffb208";
		wait for Clk_period;
		Addr <=  "0100000010111";
		Trees_din <= x"aaff8504";
		wait for Clk_period;
		Addr <=  "0100000011000";
		Trees_din <= x"005821dd";
		wait for Clk_period;
		Addr <=  "0100000011001";
		Trees_din <= x"ffba21dd";
		wait for Clk_period;
		Addr <=  "0100000011010";
		Trees_din <= x"ba003704";
		wait for Clk_period;
		Addr <=  "0100000011011";
		Trees_din <= x"ff8521dd";
		wait for Clk_period;
		Addr <=  "0100000011100";
		Trees_din <= x"006121dd";
		wait for Clk_period;
		Addr <=  "0100000011101";
		Trees_din <= x"adff2b08";
		wait for Clk_period;
		Addr <=  "0100000011110";
		Trees_din <= x"7cff9e04";
		wait for Clk_period;
		Addr <=  "0100000011111";
		Trees_din <= x"ff8c21dd";
		wait for Clk_period;
		Addr <=  "0100000100000";
		Trees_din <= x"002821dd";
		wait for Clk_period;
		Addr <=  "0100000100001";
		Trees_din <= x"2bffc404";
		wait for Clk_period;
		Addr <=  "0100000100010";
		Trees_din <= x"000821dd";
		wait for Clk_period;
		Addr <=  "0100000100011";
		Trees_din <= x"005621dd";
		wait for Clk_period;
		Addr <=  "0100000100100";
		Trees_din <= x"de006210";
		wait for Clk_period;
		Addr <=  "0100000100101";
		Trees_din <= x"1bffb808";
		wait for Clk_period;
		Addr <=  "0100000100110";
		Trees_din <= x"9effad04";
		wait for Clk_period;
		Addr <=  "0100000100111";
		Trees_din <= x"003721dd";
		wait for Clk_period;
		Addr <=  "0100000101000";
		Trees_din <= x"ffa721dd";
		wait for Clk_period;
		Addr <=  "0100000101001";
		Trees_din <= x"efffaa04";
		wait for Clk_period;
		Addr <=  "0100000101010";
		Trees_din <= x"fff221dd";
		wait for Clk_period;
		Addr <=  "0100000101011";
		Trees_din <= x"ff7b21dd";
		wait for Clk_period;
		Addr <=  "0100000101100";
		Trees_din <= x"79ff1808";
		wait for Clk_period;
		Addr <=  "0100000101101";
		Trees_din <= x"12ffab04";
		wait for Clk_period;
		Addr <=  "0100000101110";
		Trees_din <= x"008821dd";
		wait for Clk_period;
		Addr <=  "0100000101111";
		Trees_din <= x"ffac21dd";
		wait for Clk_period;
		Addr <=  "0100000110000";
		Trees_din <= x"48008804";
		wait for Clk_period;
		Addr <=  "0100000110001";
		Trees_din <= x"ff3f21dd";
		wait for Clk_period;
		Addr <=  "0100000110010";
		Trees_din <= x"002521dd";
		wait for Clk_period;
		Addr <=  "0100000110011";
		Trees_din <= x"53fffe20";
		wait for Clk_period;
		Addr <=  "0100000110100";
		Trees_din <= x"d700dd10";
		wait for Clk_period;
		Addr <=  "0100000110101";
		Trees_din <= x"b2ffd108";
		wait for Clk_period;
		Addr <=  "0100000110110";
		Trees_din <= x"9bffee04";
		wait for Clk_period;
		Addr <=  "0100000110111";
		Trees_din <= x"001c21dd";
		wait for Clk_period;
		Addr <=  "0100000111000";
		Trees_din <= x"ffb321dd";
		wait for Clk_period;
		Addr <=  "0100000111001";
		Trees_din <= x"7dfff504";
		wait for Clk_period;
		Addr <=  "0100000111010";
		Trees_din <= x"005021dd";
		wait for Clk_period;
		Addr <=  "0100000111011";
		Trees_din <= x"000121dd";
		wait for Clk_period;
		Addr <=  "0100000111100";
		Trees_din <= x"dfff7408";
		wait for Clk_period;
		Addr <=  "0100000111101";
		Trees_din <= x"b0ff3f04";
		wait for Clk_period;
		Addr <=  "0100000111110";
		Trees_din <= x"007321dd";
		wait for Clk_period;
		Addr <=  "0100000111111";
		Trees_din <= x"ff9a21dd";
		wait for Clk_period;
		Addr <=  "0100001000000";
		Trees_din <= x"81ffba04";
		wait for Clk_period;
		Addr <=  "0100001000001";
		Trees_din <= x"ff6621dd";
		wait for Clk_period;
		Addr <=  "0100001000010";
		Trees_din <= x"000b21dd";
		wait for Clk_period;
		Addr <=  "0100001000011";
		Trees_din <= x"4cffa610";
		wait for Clk_period;
		Addr <=  "0100001000100";
		Trees_din <= x"26001f08";
		wait for Clk_period;
		Addr <=  "0100001000101";
		Trees_din <= x"e1003b04";
		wait for Clk_period;
		Addr <=  "0100001000110";
		Trees_din <= x"009921dd";
		wait for Clk_period;
		Addr <=  "0100001000111";
		Trees_din <= x"ffc421dd";
		wait for Clk_period;
		Addr <=  "0100001001000";
		Trees_din <= x"1cffa804";
		wait for Clk_period;
		Addr <=  "0100001001001";
		Trees_din <= x"ff9921dd";
		wait for Clk_period;
		Addr <=  "0100001001010";
		Trees_din <= x"003421dd";
		wait for Clk_period;
		Addr <=  "0100001001011";
		Trees_din <= x"ff5c21dd";
		wait for Clk_period;
		Addr <=  "0100001001100";
		Trees_din <= x"da007b40";
		wait for Clk_period;
		Addr <=  "0100001001101";
		Trees_din <= x"e5fee420";
		wait for Clk_period;
		Addr <=  "0100001001110";
		Trees_din <= x"a8ffb710";
		wait for Clk_period;
		Addr <=  "0100001001111";
		Trees_din <= x"50ff7208";
		wait for Clk_period;
		Addr <=  "0100001010000";
		Trees_din <= x"05001504";
		wait for Clk_period;
		Addr <=  "0100001010001";
		Trees_din <= x"001621dd";
		wait for Clk_period;
		Addr <=  "0100001010010";
		Trees_din <= x"ffa021dd";
		wait for Clk_period;
		Addr <=  "0100001010011";
		Trees_din <= x"98ff3a04";
		wait for Clk_period;
		Addr <=  "0100001010100";
		Trees_din <= x"ffd421dd";
		wait for Clk_period;
		Addr <=  "0100001010101";
		Trees_din <= x"003621dd";
		wait for Clk_period;
		Addr <=  "0100001010110";
		Trees_din <= x"01fea808";
		wait for Clk_period;
		Addr <=  "0100001010111";
		Trees_din <= x"74003304";
		wait for Clk_period;
		Addr <=  "0100001011000";
		Trees_din <= x"ffa821dd";
		wait for Clk_period;
		Addr <=  "0100001011001";
		Trees_din <= x"006e21dd";
		wait for Clk_period;
		Addr <=  "0100001011010";
		Trees_din <= x"e7001204";
		wait for Clk_period;
		Addr <=  "0100001011011";
		Trees_din <= x"006721dd";
		wait for Clk_period;
		Addr <=  "0100001011100";
		Trees_din <= x"ff9921dd";
		wait for Clk_period;
		Addr <=  "0100001011101";
		Trees_din <= x"4effb710";
		wait for Clk_period;
		Addr <=  "0100001011110";
		Trees_din <= x"f8006a08";
		wait for Clk_period;
		Addr <=  "0100001011111";
		Trees_din <= x"c2ffc604";
		wait for Clk_period;
		Addr <=  "0100001100000";
		Trees_din <= x"002621dd";
		wait for Clk_period;
		Addr <=  "0100001100001";
		Trees_din <= x"ff9521dd";
		wait for Clk_period;
		Addr <=  "0100001100010";
		Trees_din <= x"9dff2204";
		wait for Clk_period;
		Addr <=  "0100001100011";
		Trees_din <= x"ffd921dd";
		wait for Clk_period;
		Addr <=  "0100001100100";
		Trees_din <= x"006e21dd";
		wait for Clk_period;
		Addr <=  "0100001100101";
		Trees_din <= x"d7006708";
		wait for Clk_period;
		Addr <=  "0100001100110";
		Trees_din <= x"63ffde04";
		wait for Clk_period;
		Addr <=  "0100001100111";
		Trees_din <= x"003321dd";
		wait for Clk_period;
		Addr <=  "0100001101000";
		Trees_din <= x"ff8421dd";
		wait for Clk_period;
		Addr <=  "0100001101001";
		Trees_din <= x"d700a204";
		wait for Clk_period;
		Addr <=  "0100001101010";
		Trees_din <= x"ff5721dd";
		wait for Clk_period;
		Addr <=  "0100001101011";
		Trees_din <= x"ffce21dd";
		wait for Clk_period;
		Addr <=  "0100001101100";
		Trees_din <= x"e2ff6510";
		wait for Clk_period;
		Addr <=  "0100001101101";
		Trees_din <= x"d6001c08";
		wait for Clk_period;
		Addr <=  "0100001101110";
		Trees_din <= x"8effdc04";
		wait for Clk_period;
		Addr <=  "0100001101111";
		Trees_din <= x"ffa421dd";
		wait for Clk_period;
		Addr <=  "0100001110000";
		Trees_din <= x"006121dd";
		wait for Clk_period;
		Addr <=  "0100001110001";
		Trees_din <= x"4bfe8604";
		wait for Clk_period;
		Addr <=  "0100001110010";
		Trees_din <= x"ffe521dd";
		wait for Clk_period;
		Addr <=  "0100001110011";
		Trees_din <= x"ff4721dd";
		wait for Clk_period;
		Addr <=  "0100001110100";
		Trees_din <= x"edffcf04";
		wait for Clk_period;
		Addr <=  "0100001110101";
		Trees_din <= x"005621dd";
		wait for Clk_period;
		Addr <=  "0100001110110";
		Trees_din <= x"ffb221dd";
		wait for Clk_period;
		Addr <=  "0100001110111";
		Trees_din <= x"3100b680";
		wait for Clk_period;
		Addr <=  "0100001111000";
		Trees_din <= x"63ffd240";
		wait for Clk_period;
		Addr <=  "0100001111001";
		Trees_din <= x"3fffb420";
		wait for Clk_period;
		Addr <=  "0100001111010";
		Trees_din <= x"e7ff3010";
		wait for Clk_period;
		Addr <=  "0100001111011";
		Trees_din <= x"25001b08";
		wait for Clk_period;
		Addr <=  "0100001111100";
		Trees_din <= x"4dfe5504";
		wait for Clk_period;
		Addr <=  "0100001111101";
		Trees_din <= x"ffa82339";
		wait for Clk_period;
		Addr <=  "0100001111110";
		Trees_din <= x"007b2339";
		wait for Clk_period;
		Addr <=  "0100001111111";
		Trees_din <= x"74ffb904";
		wait for Clk_period;
		Addr <=  "0100010000000";
		Trees_din <= x"00092339";
		wait for Clk_period;
		Addr <=  "0100010000001";
		Trees_din <= x"ff4d2339";
		wait for Clk_period;
		Addr <=  "0100010000010";
		Trees_din <= x"9dff9108";
		wait for Clk_period;
		Addr <=  "0100010000011";
		Trees_din <= x"4cffb504";
		wait for Clk_period;
		Addr <=  "0100010000100";
		Trees_din <= x"00832339";
		wait for Clk_period;
		Addr <=  "0100010000101";
		Trees_din <= x"ffb02339";
		wait for Clk_period;
		Addr <=  "0100010000110";
		Trees_din <= x"06ff5504";
		wait for Clk_period;
		Addr <=  "0100010000111";
		Trees_din <= x"ffc92339";
		wait for Clk_period;
		Addr <=  "0100010001000";
		Trees_din <= x"004a2339";
		wait for Clk_period;
		Addr <=  "0100010001001";
		Trees_din <= x"5900a710";
		wait for Clk_period;
		Addr <=  "0100010001010";
		Trees_din <= x"b4ff6e08";
		wait for Clk_period;
		Addr <=  "0100010001011";
		Trees_din <= x"0cff4604";
		wait for Clk_period;
		Addr <=  "0100010001100";
		Trees_din <= x"ffff2339";
		wait for Clk_period;
		Addr <=  "0100010001101";
		Trees_din <= x"ffbc2339";
		wait for Clk_period;
		Addr <=  "0100010001110";
		Trees_din <= x"faff9004";
		wait for Clk_period;
		Addr <=  "0100010001111";
		Trees_din <= x"00072339";
		wait for Clk_period;
		Addr <=  "0100010010000";
		Trees_din <= x"00532339";
		wait for Clk_period;
		Addr <=  "0100010010001";
		Trees_din <= x"26008e08";
		wait for Clk_period;
		Addr <=  "0100010010010";
		Trees_din <= x"9cffd904";
		wait for Clk_period;
		Addr <=  "0100010010011";
		Trees_din <= x"009a2339";
		wait for Clk_period;
		Addr <=  "0100010010100";
		Trees_din <= x"ffaa2339";
		wait for Clk_period;
		Addr <=  "0100010010101";
		Trees_din <= x"4ffec804";
		wait for Clk_period;
		Addr <=  "0100010010110";
		Trees_din <= x"004a2339";
		wait for Clk_period;
		Addr <=  "0100010010111";
		Trees_din <= x"ff6f2339";
		wait for Clk_period;
		Addr <=  "0100010011000";
		Trees_din <= x"1eff9120";
		wait for Clk_period;
		Addr <=  "0100010011001";
		Trees_din <= x"6affe210";
		wait for Clk_period;
		Addr <=  "0100010011010";
		Trees_din <= x"deffa408";
		wait for Clk_period;
		Addr <=  "0100010011011";
		Trees_din <= x"15ff0d04";
		wait for Clk_period;
		Addr <=  "0100010011100";
		Trees_din <= x"00112339";
		wait for Clk_period;
		Addr <=  "0100010011101";
		Trees_din <= x"ff642339";
		wait for Clk_period;
		Addr <=  "0100010011110";
		Trees_din <= x"36ffac04";
		wait for Clk_period;
		Addr <=  "0100010011111";
		Trees_din <= x"00232339";
		wait for Clk_period;
		Addr <=  "0100010100000";
		Trees_din <= x"ffa12339";
		wait for Clk_period;
		Addr <=  "0100010100001";
		Trees_din <= x"66ff4108";
		wait for Clk_period;
		Addr <=  "0100010100010";
		Trees_din <= x"31ff2004";
		wait for Clk_period;
		Addr <=  "0100010100011";
		Trees_din <= x"ffc12339";
		wait for Clk_period;
		Addr <=  "0100010100100";
		Trees_din <= x"00862339";
		wait for Clk_period;
		Addr <=  "0100010100101";
		Trees_din <= x"c9ff4704";
		wait for Clk_period;
		Addr <=  "0100010100110";
		Trees_din <= x"00032339";
		wait for Clk_period;
		Addr <=  "0100010100111";
		Trees_din <= x"ff652339";
		wait for Clk_period;
		Addr <=  "0100010101000";
		Trees_din <= x"09ffe910";
		wait for Clk_period;
		Addr <=  "0100010101001";
		Trees_din <= x"b7ffb508";
		wait for Clk_period;
		Addr <=  "0100010101010";
		Trees_din <= x"1dff5a04";
		wait for Clk_period;
		Addr <=  "0100010101011";
		Trees_din <= x"00172339";
		wait for Clk_period;
		Addr <=  "0100010101100";
		Trees_din <= x"ff922339";
		wait for Clk_period;
		Addr <=  "0100010101101";
		Trees_din <= x"f8008d04";
		wait for Clk_period;
		Addr <=  "0100010101110";
		Trees_din <= x"006a2339";
		wait for Clk_period;
		Addr <=  "0100010101111";
		Trees_din <= x"ffe02339";
		wait for Clk_period;
		Addr <=  "0100010110000";
		Trees_din <= x"6e001508";
		wait for Clk_period;
		Addr <=  "0100010110001";
		Trees_din <= x"b7ff9f04";
		wait for Clk_period;
		Addr <=  "0100010110010";
		Trees_din <= x"00682339";
		wait for Clk_period;
		Addr <=  "0100010110011";
		Trees_din <= x"ffc92339";
		wait for Clk_period;
		Addr <=  "0100010110100";
		Trees_din <= x"4ffecb04";
		wait for Clk_period;
		Addr <=  "0100010110101";
		Trees_din <= x"00552339";
		wait for Clk_period;
		Addr <=  "0100010110110";
		Trees_din <= x"ff662339";
		wait for Clk_period;
		Addr <=  "0100010110111";
		Trees_din <= x"4bfe3008";
		wait for Clk_period;
		Addr <=  "0100010111000";
		Trees_din <= x"33ff4604";
		wait for Clk_period;
		Addr <=  "0100010111001";
		Trees_din <= x"000c2339";
		wait for Clk_period;
		Addr <=  "0100010111010";
		Trees_din <= x"00782339";
		wait for Clk_period;
		Addr <=  "0100010111011";
		Trees_din <= x"cffff810";
		wait for Clk_period;
		Addr <=  "0100010111100";
		Trees_din <= x"c8ffc108";
		wait for Clk_period;
		Addr <=  "0100010111101";
		Trees_din <= x"b3ff3504";
		wait for Clk_period;
		Addr <=  "0100010111110";
		Trees_din <= x"007f2339";
		wait for Clk_period;
		Addr <=  "0100010111111";
		Trees_din <= x"ffe72339";
		wait for Clk_period;
		Addr <=  "0100011000000";
		Trees_din <= x"5dffc604";
		wait for Clk_period;
		Addr <=  "0100011000001";
		Trees_din <= x"ff8a2339";
		wait for Clk_period;
		Addr <=  "0100011000010";
		Trees_din <= x"fffc2339";
		wait for Clk_period;
		Addr <=  "0100011000011";
		Trees_din <= x"37ffbd0c";
		wait for Clk_period;
		Addr <=  "0100011000100";
		Trees_din <= x"02ff5008";
		wait for Clk_period;
		Addr <=  "0100011000101";
		Trees_din <= x"40ffb804";
		wait for Clk_period;
		Addr <=  "0100011000110";
		Trees_din <= x"ffdc2339";
		wait for Clk_period;
		Addr <=  "0100011000111";
		Trees_din <= x"ff572339";
		wait for Clk_period;
		Addr <=  "0100011001000";
		Trees_din <= x"00162339";
		wait for Clk_period;
		Addr <=  "0100011001001";
		Trees_din <= x"f9ff3708";
		wait for Clk_period;
		Addr <=  "0100011001010";
		Trees_din <= x"c6ff2d04";
		wait for Clk_period;
		Addr <=  "0100011001011";
		Trees_din <= x"fff92339";
		wait for Clk_period;
		Addr <=  "0100011001100";
		Trees_din <= x"ff852339";
		wait for Clk_period;
		Addr <=  "0100011001101";
		Trees_din <= x"00652339";
		wait for Clk_period;
		Addr <=  "0100011001110";
		Trees_din <= x"31feff48";
		wait for Clk_period;
		Addr <=  "0100011001111";
		Trees_din <= x"7d004538";
		wait for Clk_period;
		Addr <=  "0100011010000";
		Trees_din <= x"20ff6c20";
		wait for Clk_period;
		Addr <=  "0100011010001";
		Trees_din <= x"bffefd10";
		wait for Clk_period;
		Addr <=  "0100011010010";
		Trees_din <= x"b9ff1408";
		wait for Clk_period;
		Addr <=  "0100011010011";
		Trees_din <= x"63ff4e04";
		wait for Clk_period;
		Addr <=  "0100011010100";
		Trees_din <= x"ffdd24bd";
		wait for Clk_period;
		Addr <=  "0100011010101";
		Trees_din <= x"008124bd";
		wait for Clk_period;
		Addr <=  "0100011010110";
		Trees_din <= x"f3fecf04";
		wait for Clk_period;
		Addr <=  "0100011010111";
		Trees_din <= x"ff6124bd";
		wait for Clk_period;
		Addr <=  "0100011011000";
		Trees_din <= x"001124bd";
		wait for Clk_period;
		Addr <=  "0100011011001";
		Trees_din <= x"2c000c08";
		wait for Clk_period;
		Addr <=  "0100011011010";
		Trees_din <= x"fafe8f04";
		wait for Clk_period;
		Addr <=  "0100011011011";
		Trees_din <= x"ffc024bd";
		wait for Clk_period;
		Addr <=  "0100011011100";
		Trees_din <= x"008524bd";
		wait for Clk_period;
		Addr <=  "0100011011101";
		Trees_din <= x"07ffce04";
		wait for Clk_period;
		Addr <=  "0100011011110";
		Trees_din <= x"005b24bd";
		wait for Clk_period;
		Addr <=  "0100011011111";
		Trees_din <= x"ff8824bd";
		wait for Clk_period;
		Addr <=  "0100011100000";
		Trees_din <= x"fbffd50c";
		wait for Clk_period;
		Addr <=  "0100011100001";
		Trees_din <= x"d0fff704";
		wait for Clk_period;
		Addr <=  "0100011100010";
		Trees_din <= x"ffa024bd";
		wait for Clk_period;
		Addr <=  "0100011100011";
		Trees_din <= x"45feb104";
		wait for Clk_period;
		Addr <=  "0100011100100";
		Trees_din <= x"ffe824bd";
		wait for Clk_period;
		Addr <=  "0100011100101";
		Trees_din <= x"009224bd";
		wait for Clk_period;
		Addr <=  "0100011100110";
		Trees_din <= x"edff6304";
		wait for Clk_period;
		Addr <=  "0100011100111";
		Trees_din <= x"006c24bd";
		wait for Clk_period;
		Addr <=  "0100011101000";
		Trees_din <= x"97ff5704";
		wait for Clk_period;
		Addr <=  "0100011101001";
		Trees_din <= x"ff7624bd";
		wait for Clk_period;
		Addr <=  "0100011101010";
		Trees_din <= x"004024bd";
		wait for Clk_period;
		Addr <=  "0100011101011";
		Trees_din <= x"8e003508";
		wait for Clk_period;
		Addr <=  "0100011101100";
		Trees_din <= x"a6ffa004";
		wait for Clk_period;
		Addr <=  "0100011101101";
		Trees_din <= x"ff6424bd";
		wait for Clk_period;
		Addr <=  "0100011101110";
		Trees_din <= x"000224bd";
		wait for Clk_period;
		Addr <=  "0100011101111";
		Trees_din <= x"5effe404";
		wait for Clk_period;
		Addr <=  "0100011110000";
		Trees_din <= x"ffe824bd";
		wait for Clk_period;
		Addr <=  "0100011110001";
		Trees_din <= x"005b24bd";
		wait for Clk_period;
		Addr <=  "0100011110010";
		Trees_din <= x"44005b40";
		wait for Clk_period;
		Addr <=  "0100011110011";
		Trees_din <= x"62ff4620";
		wait for Clk_period;
		Addr <=  "0100011110100";
		Trees_din <= x"5fffc210";
		wait for Clk_period;
		Addr <=  "0100011110101";
		Trees_din <= x"71000d08";
		wait for Clk_period;
		Addr <=  "0100011110110";
		Trees_din <= x"90ff5704";
		wait for Clk_period;
		Addr <=  "0100011110111";
		Trees_din <= x"000824bd";
		wait for Clk_period;
		Addr <=  "0100011111000";
		Trees_din <= x"ffdd24bd";
		wait for Clk_period;
		Addr <=  "0100011111001";
		Trees_din <= x"25fefc04";
		wait for Clk_period;
		Addr <=  "0100011111010";
		Trees_din <= x"003924bd";
		wait for Clk_period;
		Addr <=  "0100011111011";
		Trees_din <= x"ff6d24bd";
		wait for Clk_period;
		Addr <=  "0100011111100";
		Trees_din <= x"d1ff3508";
		wait for Clk_period;
		Addr <=  "0100011111101";
		Trees_din <= x"c8000804";
		wait for Clk_period;
		Addr <=  "0100011111110";
		Trees_din <= x"006924bd";
		wait for Clk_period;
		Addr <=  "0100011111111";
		Trees_din <= x"ffc324bd";
		wait for Clk_period;
		Addr <=  "0100100000000";
		Trees_din <= x"9dfffc04";
		wait for Clk_period;
		Addr <=  "0100100000001";
		Trees_din <= x"009024bd";
		wait for Clk_period;
		Addr <=  "0100100000010";
		Trees_din <= x"fffe24bd";
		wait for Clk_period;
		Addr <=  "0100100000011";
		Trees_din <= x"72001610";
		wait for Clk_period;
		Addr <=  "0100100000100";
		Trees_din <= x"5400fb08";
		wait for Clk_period;
		Addr <=  "0100100000101";
		Trees_din <= x"81ff9f04";
		wait for Clk_period;
		Addr <=  "0100100000110";
		Trees_din <= x"ffeb24bd";
		wait for Clk_period;
		Addr <=  "0100100000111";
		Trees_din <= x"001d24bd";
		wait for Clk_period;
		Addr <=  "0100100001000";
		Trees_din <= x"43ffa404";
		wait for Clk_period;
		Addr <=  "0100100001001";
		Trees_din <= x"ff3f24bd";
		wait for Clk_period;
		Addr <=  "0100100001010";
		Trees_din <= x"002524bd";
		wait for Clk_period;
		Addr <=  "0100100001011";
		Trees_din <= x"2fff6808";
		wait for Clk_period;
		Addr <=  "0100100001100";
		Trees_din <= x"fdfeec04";
		wait for Clk_period;
		Addr <=  "0100100001101";
		Trees_din <= x"ffe424bd";
		wait for Clk_period;
		Addr <=  "0100100001110";
		Trees_din <= x"006824bd";
		wait for Clk_period;
		Addr <=  "0100100001111";
		Trees_din <= x"2a00c904";
		wait for Clk_period;
		Addr <=  "0100100010000";
		Trees_din <= x"002524bd";
		wait for Clk_period;
		Addr <=  "0100100010001";
		Trees_din <= x"ffab24bd";
		wait for Clk_period;
		Addr <=  "0100100010010";
		Trees_din <= x"7dff7e1c";
		wait for Clk_period;
		Addr <=  "0100100010011";
		Trees_din <= x"c1fec70c";
		wait for Clk_period;
		Addr <=  "0100100010100";
		Trees_din <= x"50ff0204";
		wait for Clk_period;
		Addr <=  "0100100010101";
		Trees_din <= x"ff9124bd";
		wait for Clk_period;
		Addr <=  "0100100010110";
		Trees_din <= x"2500a504";
		wait for Clk_period;
		Addr <=  "0100100010111";
		Trees_din <= x"009824bd";
		wait for Clk_period;
		Addr <=  "0100100011000";
		Trees_din <= x"ffa124bd";
		wait for Clk_period;
		Addr <=  "0100100011001";
		Trees_din <= x"a2ffbd08";
		wait for Clk_period;
		Addr <=  "0100100011010";
		Trees_din <= x"3affbf04";
		wait for Clk_period;
		Addr <=  "0100100011011";
		Trees_din <= x"007324bd";
		wait for Clk_period;
		Addr <=  "0100100011100";
		Trees_din <= x"ffaa24bd";
		wait for Clk_period;
		Addr <=  "0100100011101";
		Trees_din <= x"a6ff3104";
		wait for Clk_period;
		Addr <=  "0100100011110";
		Trees_din <= x"002324bd";
		wait for Clk_period;
		Addr <=  "0100100011111";
		Trees_din <= x"ff4d24bd";
		wait for Clk_period;
		Addr <=  "0100100100000";
		Trees_din <= x"00fef810";
		wait for Clk_period;
		Addr <=  "0100100100001";
		Trees_din <= x"49000608";
		wait for Clk_period;
		Addr <=  "0100100100010";
		Trees_din <= x"50ff6604";
		wait for Clk_period;
		Addr <=  "0100100100011";
		Trees_din <= x"ff8224bd";
		wait for Clk_period;
		Addr <=  "0100100100100";
		Trees_din <= x"000124bd";
		wait for Clk_period;
		Addr <=  "0100100100101";
		Trees_din <= x"cf006504";
		wait for Clk_period;
		Addr <=  "0100100100110";
		Trees_din <= x"00a224bd";
		wait for Clk_period;
		Addr <=  "0100100100111";
		Trees_din <= x"ffd824bd";
		wait for Clk_period;
		Addr <=  "0100100101000";
		Trees_din <= x"66ff7408";
		wait for Clk_period;
		Addr <=  "0100100101001";
		Trees_din <= x"b7ff8504";
		wait for Clk_period;
		Addr <=  "0100100101010";
		Trees_din <= x"ff7624bd";
		wait for Clk_period;
		Addr <=  "0100100101011";
		Trees_din <= x"005024bd";
		wait for Clk_period;
		Addr <=  "0100100101100";
		Trees_din <= x"4cfede04";
		wait for Clk_period;
		Addr <=  "0100100101101";
		Trees_din <= x"fff524bd";
		wait for Clk_period;
		Addr <=  "0100100101110";
		Trees_din <= x"ff8224bd";
		wait for Clk_period;
		Addr <=  "0100100101111";
		Trees_din <= x"f5007e78";
		wait for Clk_period;
		Addr <=  "0100100110000";
		Trees_din <= x"5bff9140";
		wait for Clk_period;
		Addr <=  "0100100110001";
		Trees_din <= x"05ffea20";
		wait for Clk_period;
		Addr <=  "0100100110010";
		Trees_din <= x"4fff3a10";
		wait for Clk_period;
		Addr <=  "0100100110011";
		Trees_din <= x"c5ff5c08";
		wait for Clk_period;
		Addr <=  "0100100110100";
		Trees_din <= x"93fff204";
		wait for Clk_period;
		Addr <=  "0100100110101";
		Trees_din <= x"009325f1";
		wait for Clk_period;
		Addr <=  "0100100110110";
		Trees_din <= x"ffd025f1";
		wait for Clk_period;
		Addr <=  "0100100110111";
		Trees_din <= x"b1ff1a04";
		wait for Clk_period;
		Addr <=  "0100100111000";
		Trees_din <= x"ff9925f1";
		wait for Clk_period;
		Addr <=  "0100100111001";
		Trees_din <= x"005d25f1";
		wait for Clk_period;
		Addr <=  "0100100111010";
		Trees_din <= x"00ff4b08";
		wait for Clk_period;
		Addr <=  "0100100111011";
		Trees_din <= x"7d001604";
		wait for Clk_period;
		Addr <=  "0100100111100";
		Trees_din <= x"006425f1";
		wait for Clk_period;
		Addr <=  "0100100111101";
		Trees_din <= x"ff9b25f1";
		wait for Clk_period;
		Addr <=  "0100100111110";
		Trees_din <= x"2dfe9204";
		wait for Clk_period;
		Addr <=  "0100100111111";
		Trees_din <= x"ff7025f1";
		wait for Clk_period;
		Addr <=  "0100101000000";
		Trees_din <= x"fffe25f1";
		wait for Clk_period;
		Addr <=  "0100101000001";
		Trees_din <= x"91ff7510";
		wait for Clk_period;
		Addr <=  "0100101000010";
		Trees_din <= x"beffa008";
		wait for Clk_period;
		Addr <=  "0100101000011";
		Trees_din <= x"d8004304";
		wait for Clk_period;
		Addr <=  "0100101000100";
		Trees_din <= x"003425f1";
		wait for Clk_period;
		Addr <=  "0100101000101";
		Trees_din <= x"ffcc25f1";
		wait for Clk_period;
		Addr <=  "0100101000110";
		Trees_din <= x"c9ff8f04";
		wait for Clk_period;
		Addr <=  "0100101000111";
		Trees_din <= x"000025f1";
		wait for Clk_period;
		Addr <=  "0100101001000";
		Trees_din <= x"ffb225f1";
		wait for Clk_period;
		Addr <=  "0100101001001";
		Trees_din <= x"3eff9a08";
		wait for Clk_period;
		Addr <=  "0100101001010";
		Trees_din <= x"fa000504";
		wait for Clk_period;
		Addr <=  "0100101001011";
		Trees_din <= x"001325f1";
		wait for Clk_period;
		Addr <=  "0100101001100";
		Trees_din <= x"ffac25f1";
		wait for Clk_period;
		Addr <=  "0100101001101";
		Trees_din <= x"57ffa604";
		wait for Clk_period;
		Addr <=  "0100101001110";
		Trees_din <= x"ffc125f1";
		wait for Clk_period;
		Addr <=  "0100101001111";
		Trees_din <= x"004e25f1";
		wait for Clk_period;
		Addr <=  "0100101010000";
		Trees_din <= x"b9ff7b1c";
		wait for Clk_period;
		Addr <=  "0100101010001";
		Trees_din <= x"32ff5310";
		wait for Clk_period;
		Addr <=  "0100101010010";
		Trees_din <= x"0cff4a08";
		wait for Clk_period;
		Addr <=  "0100101010011";
		Trees_din <= x"c2ff7304";
		wait for Clk_period;
		Addr <=  "0100101010100";
		Trees_din <= x"003125f1";
		wait for Clk_period;
		Addr <=  "0100101010101";
		Trees_din <= x"fffc25f1";
		wait for Clk_period;
		Addr <=  "0100101010110";
		Trees_din <= x"a0fe3804";
		wait for Clk_period;
		Addr <=  "0100101010111";
		Trees_din <= x"002b25f1";
		wait for Clk_period;
		Addr <=  "0100101011000";
		Trees_din <= x"ff6b25f1";
		wait for Clk_period;
		Addr <=  "0100101011001";
		Trees_din <= x"afff5804";
		wait for Clk_period;
		Addr <=  "0100101011010";
		Trees_din <= x"ffbf25f1";
		wait for Clk_period;
		Addr <=  "0100101011011";
		Trees_din <= x"50ff3704";
		wait for Clk_period;
		Addr <=  "0100101011100";
		Trees_din <= x"001825f1";
		wait for Clk_period;
		Addr <=  "0100101011101";
		Trees_din <= x"008d25f1";
		wait for Clk_period;
		Addr <=  "0100101011110";
		Trees_din <= x"37fff810";
		wait for Clk_period;
		Addr <=  "0100101011111";
		Trees_din <= x"e1fffe08";
		wait for Clk_period;
		Addr <=  "0100101100000";
		Trees_din <= x"2fff4904";
		wait for Clk_period;
		Addr <=  "0100101100001";
		Trees_din <= x"002525f1";
		wait for Clk_period;
		Addr <=  "0100101100010";
		Trees_din <= x"ff7b25f1";
		wait for Clk_period;
		Addr <=  "0100101100011";
		Trees_din <= x"a3ffdc04";
		wait for Clk_period;
		Addr <=  "0100101100100";
		Trees_din <= x"006025f1";
		wait for Clk_period;
		Addr <=  "0100101100101";
		Trees_din <= x"ff8b25f1";
		wait for Clk_period;
		Addr <=  "0100101100110";
		Trees_din <= x"62ffc408";
		wait for Clk_period;
		Addr <=  "0100101100111";
		Trees_din <= x"1cffdc04";
		wait for Clk_period;
		Addr <=  "0100101101000";
		Trees_din <= x"008625f1";
		wait for Clk_period;
		Addr <=  "0100101101001";
		Trees_din <= x"ffd825f1";
		wait for Clk_period;
		Addr <=  "0100101101010";
		Trees_din <= x"ff9225f1";
		wait for Clk_period;
		Addr <=  "0100101101011";
		Trees_din <= x"2dff4318";
		wait for Clk_period;
		Addr <=  "0100101101100";
		Trees_din <= x"bf000f10";
		wait for Clk_period;
		Addr <=  "0100101101101";
		Trees_din <= x"ee00c40c";
		wait for Clk_period;
		Addr <=  "0100101101110";
		Trees_din <= x"20008708";
		wait for Clk_period;
		Addr <=  "0100101101111";
		Trees_din <= x"05ffce04";
		wait for Clk_period;
		Addr <=  "0100101110000";
		Trees_din <= x"ffe025f1";
		wait for Clk_period;
		Addr <=  "0100101110001";
		Trees_din <= x"008e25f1";
		wait for Clk_period;
		Addr <=  "0100101110010";
		Trees_din <= x"ffd125f1";
		wait for Clk_period;
		Addr <=  "0100101110011";
		Trees_din <= x"ffb525f1";
		wait for Clk_period;
		Addr <=  "0100101110100";
		Trees_din <= x"c8fffa04";
		wait for Clk_period;
		Addr <=  "0100101110101";
		Trees_din <= x"002c25f1";
		wait for Clk_period;
		Addr <=  "0100101110110";
		Trees_din <= x"ff7c25f1";
		wait for Clk_period;
		Addr <=  "0100101110111";
		Trees_din <= x"77fede04";
		wait for Clk_period;
		Addr <=  "0100101111000";
		Trees_din <= x"001f25f1";
		wait for Clk_period;
		Addr <=  "0100101111001";
		Trees_din <= x"cf001f04";
		wait for Clk_period;
		Addr <=  "0100101111010";
		Trees_din <= x"ffeb25f1";
		wait for Clk_period;
		Addr <=  "0100101111011";
		Trees_din <= x"ff8525f1";
		wait for Clk_period;
		Addr <=  "0100101111100";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0100101111101";
		Trees_din <= x"40005868";
		wait for Clk_period;
		Addr <=  "0100101111110";
		Trees_din <= x"cafdaa28";
		wait for Clk_period;
		Addr <=  "0100101111111";
		Trees_din <= x"17007720";
		wait for Clk_period;
		Addr <=  "0100110000000";
		Trees_din <= x"37ffe410";
		wait for Clk_period;
		Addr <=  "0100110000001";
		Trees_din <= x"b0ffdb08";
		wait for Clk_period;
		Addr <=  "0100110000010";
		Trees_din <= x"60ff0b04";
		wait for Clk_period;
		Addr <=  "0100110000011";
		Trees_din <= x"00392741";
		wait for Clk_period;
		Addr <=  "0100110000100";
		Trees_din <= x"ff7b2741";
		wait for Clk_period;
		Addr <=  "0100110000101";
		Trees_din <= x"69ff2f04";
		wait for Clk_period;
		Addr <=  "0100110000110";
		Trees_din <= x"ffb92741";
		wait for Clk_period;
		Addr <=  "0100110000111";
		Trees_din <= x"006f2741";
		wait for Clk_period;
		Addr <=  "0100110001000";
		Trees_din <= x"99fe1808";
		wait for Clk_period;
		Addr <=  "0100110001001";
		Trees_din <= x"fcff0904";
		wait for Clk_period;
		Addr <=  "0100110001010";
		Trees_din <= x"ff742741";
		wait for Clk_period;
		Addr <=  "0100110001011";
		Trees_din <= x"fff62741";
		wait for Clk_period;
		Addr <=  "0100110001100";
		Trees_din <= x"41fecb04";
		wait for Clk_period;
		Addr <=  "0100110001101";
		Trees_din <= x"007e2741";
		wait for Clk_period;
		Addr <=  "0100110001110";
		Trees_din <= x"ffe42741";
		wait for Clk_period;
		Addr <=  "0100110001111";
		Trees_din <= x"24ff4d04";
		wait for Clk_period;
		Addr <=  "0100110010000";
		Trees_din <= x"ffcb2741";
		wait for Clk_period;
		Addr <=  "0100110010001";
		Trees_din <= x"008e2741";
		wait for Clk_period;
		Addr <=  "0100110010010";
		Trees_din <= x"9bff3b20";
		wait for Clk_period;
		Addr <=  "0100110010011";
		Trees_din <= x"17fffe10";
		wait for Clk_period;
		Addr <=  "0100110010100";
		Trees_din <= x"a5ff3608";
		wait for Clk_period;
		Addr <=  "0100110010101";
		Trees_din <= x"94ffcf04";
		wait for Clk_period;
		Addr <=  "0100110010110";
		Trees_din <= x"ffb32741";
		wait for Clk_period;
		Addr <=  "0100110010111";
		Trees_din <= x"fffb2741";
		wait for Clk_period;
		Addr <=  "0100110011000";
		Trees_din <= x"a1ffc804";
		wait for Clk_period;
		Addr <=  "0100110011001";
		Trees_din <= x"002e2741";
		wait for Clk_period;
		Addr <=  "0100110011010";
		Trees_din <= x"ff942741";
		wait for Clk_period;
		Addr <=  "0100110011011";
		Trees_din <= x"21ffc808";
		wait for Clk_period;
		Addr <=  "0100110011100";
		Trees_din <= x"25009404";
		wait for Clk_period;
		Addr <=  "0100110011101";
		Trees_din <= x"00022741";
		wait for Clk_period;
		Addr <=  "0100110011110";
		Trees_din <= x"ff782741";
		wait for Clk_period;
		Addr <=  "0100110011111";
		Trees_din <= x"b5fece04";
		wait for Clk_period;
		Addr <=  "0100110100000";
		Trees_din <= x"00022741";
		wait for Clk_period;
		Addr <=  "0100110100001";
		Trees_din <= x"00572741";
		wait for Clk_period;
		Addr <=  "0100110100010";
		Trees_din <= x"bcff6110";
		wait for Clk_period;
		Addr <=  "0100110100011";
		Trees_din <= x"69feb908";
		wait for Clk_period;
		Addr <=  "0100110100100";
		Trees_din <= x"09fe8c04";
		wait for Clk_period;
		Addr <=  "0100110100101";
		Trees_din <= x"00522741";
		wait for Clk_period;
		Addr <=  "0100110100110";
		Trees_din <= x"ff912741";
		wait for Clk_period;
		Addr <=  "0100110100111";
		Trees_din <= x"a5ff0204";
		wait for Clk_period;
		Addr <=  "0100110101000";
		Trees_din <= x"fffc2741";
		wait for Clk_period;
		Addr <=  "0100110101001";
		Trees_din <= x"00262741";
		wait for Clk_period;
		Addr <=  "0100110101010";
		Trees_din <= x"cafeea08";
		wait for Clk_period;
		Addr <=  "0100110101011";
		Trees_din <= x"fafeb904";
		wait for Clk_period;
		Addr <=  "0100110101100";
		Trees_din <= x"ffb12741";
		wait for Clk_period;
		Addr <=  "0100110101101";
		Trees_din <= x"00492741";
		wait for Clk_period;
		Addr <=  "0100110101110";
		Trees_din <= x"5bff3004";
		wait for Clk_period;
		Addr <=  "0100110101111";
		Trees_din <= x"ff892741";
		wait for Clk_period;
		Addr <=  "0100110110000";
		Trees_din <= x"00172741";
		wait for Clk_period;
		Addr <=  "0100110110001";
		Trees_din <= x"1aff141c";
		wait for Clk_period;
		Addr <=  "0100110110010";
		Trees_din <= x"65fff514";
		wait for Clk_period;
		Addr <=  "0100110110011";
		Trees_din <= x"4800a110";
		wait for Clk_period;
		Addr <=  "0100110110100";
		Trees_din <= x"77ff3008";
		wait for Clk_period;
		Addr <=  "0100110110101";
		Trees_din <= x"5ffe9304";
		wait for Clk_period;
		Addr <=  "0100110110110";
		Trees_din <= x"002d2741";
		wait for Clk_period;
		Addr <=  "0100110110111";
		Trees_din <= x"ff742741";
		wait for Clk_period;
		Addr <=  "0100110111000";
		Trees_din <= x"dc002304";
		wait for Clk_period;
		Addr <=  "0100110111001";
		Trees_din <= x"00062741";
		wait for Clk_period;
		Addr <=  "0100110111010";
		Trees_din <= x"ff8c2741";
		wait for Clk_period;
		Addr <=  "0100110111011";
		Trees_din <= x"006f2741";
		wait for Clk_period;
		Addr <=  "0100110111100";
		Trees_din <= x"feff6c04";
		wait for Clk_period;
		Addr <=  "0100110111101";
		Trees_din <= x"007a2741";
		wait for Clk_period;
		Addr <=  "0100110111110";
		Trees_din <= x"fffa2741";
		wait for Clk_period;
		Addr <=  "0100110111111";
		Trees_din <= x"48ff7e0c";
		wait for Clk_period;
		Addr <=  "0100111000000";
		Trees_din <= x"8b003108";
		wait for Clk_period;
		Addr <=  "0100111000001";
		Trees_din <= x"18000004";
		wait for Clk_period;
		Addr <=  "0100111000010";
		Trees_din <= x"ff662741";
		wait for Clk_period;
		Addr <=  "0100111000011";
		Trees_din <= x"000c2741";
		wait for Clk_period;
		Addr <=  "0100111000100";
		Trees_din <= x"00472741";
		wait for Clk_period;
		Addr <=  "0100111000101";
		Trees_din <= x"f9feae08";
		wait for Clk_period;
		Addr <=  "0100111000110";
		Trees_din <= x"0cfebf04";
		wait for Clk_period;
		Addr <=  "0100111000111";
		Trees_din <= x"ff892741";
		wait for Clk_period;
		Addr <=  "0100111001000";
		Trees_din <= x"00052741";
		wait for Clk_period;
		Addr <=  "0100111001001";
		Trees_din <= x"6bfe3108";
		wait for Clk_period;
		Addr <=  "0100111001010";
		Trees_din <= x"ecffc404";
		wait for Clk_period;
		Addr <=  "0100111001011";
		Trees_din <= x"ff832741";
		wait for Clk_period;
		Addr <=  "0100111001100";
		Trees_din <= x"00172741";
		wait for Clk_period;
		Addr <=  "0100111001101";
		Trees_din <= x"60ffc904";
		wait for Clk_period;
		Addr <=  "0100111001110";
		Trees_din <= x"00792741";
		wait for Clk_period;
		Addr <=  "0100111001111";
		Trees_din <= x"fff42741";
		wait for Clk_period;
		Addr <=  "0100111010000";
		Trees_din <= x"6700017c";
		wait for Clk_period;
		Addr <=  "0100111010001";
		Trees_din <= x"67ffa440";
		wait for Clk_period;
		Addr <=  "0100111010010";
		Trees_din <= x"5a001320";
		wait for Clk_period;
		Addr <=  "0100111010011";
		Trees_din <= x"24ffe810";
		wait for Clk_period;
		Addr <=  "0100111010100";
		Trees_din <= x"c8fff408";
		wait for Clk_period;
		Addr <=  "0100111010101";
		Trees_din <= x"bfff4004";
		wait for Clk_period;
		Addr <=  "0100111010110";
		Trees_din <= x"ff8f2885";
		wait for Clk_period;
		Addr <=  "0100111010111";
		Trees_din <= x"00182885";
		wait for Clk_period;
		Addr <=  "0100111011000";
		Trees_din <= x"faff2304";
		wait for Clk_period;
		Addr <=  "0100111011001";
		Trees_din <= x"00082885";
		wait for Clk_period;
		Addr <=  "0100111011010";
		Trees_din <= x"ff7a2885";
		wait for Clk_period;
		Addr <=  "0100111011011";
		Trees_din <= x"f7ff7108";
		wait for Clk_period;
		Addr <=  "0100111011100";
		Trees_din <= x"a7ff4804";
		wait for Clk_period;
		Addr <=  "0100111011101";
		Trees_din <= x"00612885";
		wait for Clk_period;
		Addr <=  "0100111011110";
		Trees_din <= x"ff982885";
		wait for Clk_period;
		Addr <=  "0100111011111";
		Trees_din <= x"77ff4904";
		wait for Clk_period;
		Addr <=  "0100111100000";
		Trees_din <= x"008a2885";
		wait for Clk_period;
		Addr <=  "0100111100001";
		Trees_din <= x"ffdf2885";
		wait for Clk_period;
		Addr <=  "0100111100010";
		Trees_din <= x"31006710";
		wait for Clk_period;
		Addr <=  "0100111100011";
		Trees_din <= x"29ff9808";
		wait for Clk_period;
		Addr <=  "0100111100100";
		Trees_din <= x"2dff6e04";
		wait for Clk_period;
		Addr <=  "0100111100101";
		Trees_din <= x"ffff2885";
		wait for Clk_period;
		Addr <=  "0100111100110";
		Trees_din <= x"004f2885";
		wait for Clk_period;
		Addr <=  "0100111100111";
		Trees_din <= x"ebfece04";
		wait for Clk_period;
		Addr <=  "0100111101000";
		Trees_din <= x"005e2885";
		wait for Clk_period;
		Addr <=  "0100111101001";
		Trees_din <= x"00152885";
		wait for Clk_period;
		Addr <=  "0100111101010";
		Trees_din <= x"d1ff2608";
		wait for Clk_period;
		Addr <=  "0100111101011";
		Trees_din <= x"c1fec704";
		wait for Clk_period;
		Addr <=  "0100111101100";
		Trees_din <= x"ff5e2885";
		wait for Clk_period;
		Addr <=  "0100111101101";
		Trees_din <= x"fff32885";
		wait for Clk_period;
		Addr <=  "0100111101110";
		Trees_din <= x"34fff504";
		wait for Clk_period;
		Addr <=  "0100111101111";
		Trees_din <= x"00532885";
		wait for Clk_period;
		Addr <=  "0100111110000";
		Trees_din <= x"ffd12885";
		wait for Clk_period;
		Addr <=  "0100111110001";
		Trees_din <= x"5bffcb20";
		wait for Clk_period;
		Addr <=  "0100111110010";
		Trees_din <= x"44005b10";
		wait for Clk_period;
		Addr <=  "0100111110011";
		Trees_din <= x"49fff908";
		wait for Clk_period;
		Addr <=  "0100111110100";
		Trees_din <= x"26fffd04";
		wait for Clk_period;
		Addr <=  "0100111110101";
		Trees_din <= x"00372885";
		wait for Clk_period;
		Addr <=  "0100111110110";
		Trees_din <= x"ffb72885";
		wait for Clk_period;
		Addr <=  "0100111110111";
		Trees_din <= x"0cfec104";
		wait for Clk_period;
		Addr <=  "0100111111000";
		Trees_din <= x"ffe42885";
		wait for Clk_period;
		Addr <=  "0100111111001";
		Trees_din <= x"00422885";
		wait for Clk_period;
		Addr <=  "0100111111010";
		Trees_din <= x"58ff3c08";
		wait for Clk_period;
		Addr <=  "0100111111011";
		Trees_din <= x"86fe9004";
		wait for Clk_period;
		Addr <=  "0100111111100";
		Trees_din <= x"000c2885";
		wait for Clk_period;
		Addr <=  "0100111111101";
		Trees_din <= x"ff5e2885";
		wait for Clk_period;
		Addr <=  "0100111111110";
		Trees_din <= x"feff6f04";
		wait for Clk_period;
		Addr <=  "0100111111111";
		Trees_din <= x"00752885";
		wait for Clk_period;
		Addr <=  "0101000000000";
		Trees_din <= x"ffda2885";
		wait for Clk_period;
		Addr <=  "0101000000001";
		Trees_din <= x"edff8110";
		wait for Clk_period;
		Addr <=  "0101000000010";
		Trees_din <= x"cdffe308";
		wait for Clk_period;
		Addr <=  "0101000000011";
		Trees_din <= x"d1ff2c04";
		wait for Clk_period;
		Addr <=  "0101000000100";
		Trees_din <= x"ff7b2885";
		wait for Clk_period;
		Addr <=  "0101000000101";
		Trees_din <= x"00052885";
		wait for Clk_period;
		Addr <=  "0101000000110";
		Trees_din <= x"74ffc704";
		wait for Clk_period;
		Addr <=  "0101000000111";
		Trees_din <= x"00122885";
		wait for Clk_period;
		Addr <=  "0101000001000";
		Trees_din <= x"006a2885";
		wait for Clk_period;
		Addr <=  "0101000001001";
		Trees_din <= x"f4fe7b04";
		wait for Clk_period;
		Addr <=  "0101000001010";
		Trees_din <= x"ffb82885";
		wait for Clk_period;
		Addr <=  "0101000001011";
		Trees_din <= x"a3ff3704";
		wait for Clk_period;
		Addr <=  "0101000001100";
		Trees_din <= x"00142885";
		wait for Clk_period;
		Addr <=  "0101000001101";
		Trees_din <= x"00962885";
		wait for Clk_period;
		Addr <=  "0101000001110";
		Trees_din <= x"89009924";
		wait for Clk_period;
		Addr <=  "0101000001111";
		Trees_din <= x"8bffa404";
		wait for Clk_period;
		Addr <=  "0101000010000";
		Trees_din <= x"ff842885";
		wait for Clk_period;
		Addr <=  "0101000010001";
		Trees_din <= x"fbff4c10";
		wait for Clk_period;
		Addr <=  "0101000010010";
		Trees_din <= x"8ffefa08";
		wait for Clk_period;
		Addr <=  "0101000010011";
		Trees_din <= x"a2ff8c04";
		wait for Clk_period;
		Addr <=  "0101000010100";
		Trees_din <= x"ffa12885";
		wait for Clk_period;
		Addr <=  "0101000010101";
		Trees_din <= x"005b2885";
		wait for Clk_period;
		Addr <=  "0101000010110";
		Trees_din <= x"58ff1d04";
		wait for Clk_period;
		Addr <=  "0101000010111";
		Trees_din <= x"ff672885";
		wait for Clk_period;
		Addr <=  "0101000011000";
		Trees_din <= x"000c2885";
		wait for Clk_period;
		Addr <=  "0101000011001";
		Trees_din <= x"87ff3c08";
		wait for Clk_period;
		Addr <=  "0101000011010";
		Trees_din <= x"65ff2704";
		wait for Clk_period;
		Addr <=  "0101000011011";
		Trees_din <= x"ff6f2885";
		wait for Clk_period;
		Addr <=  "0101000011100";
		Trees_din <= x"00412885";
		wait for Clk_period;
		Addr <=  "0101000011101";
		Trees_din <= x"adffde04";
		wait for Clk_period;
		Addr <=  "0101000011110";
		Trees_din <= x"00772885";
		wait for Clk_period;
		Addr <=  "0101000011111";
		Trees_din <= x"fffb2885";
		wait for Clk_period;
		Addr <=  "0101000100000";
		Trees_din <= x"ff832885";
		wait for Clk_period;
		Addr <=  "0101000100001";
		Trees_din <= x"3d003378";
		wait for Clk_period;
		Addr <=  "0101000100010";
		Trees_din <= x"ddfedf3c";
		wait for Clk_period;
		Addr <=  "0101000100011";
		Trees_din <= x"20ff5c1c";
		wait for Clk_period;
		Addr <=  "0101000100100";
		Trees_din <= x"f2037610";
		wait for Clk_period;
		Addr <=  "0101000100101";
		Trees_din <= x"ceff9e08";
		wait for Clk_period;
		Addr <=  "0101000100110";
		Trees_din <= x"3f001404";
		wait for Clk_period;
		Addr <=  "0101000100111";
		Trees_din <= x"00512a19";
		wait for Clk_period;
		Addr <=  "0101000101000";
		Trees_din <= x"ffe22a19";
		wait for Clk_period;
		Addr <=  "0101000101001";
		Trees_din <= x"09fee604";
		wait for Clk_period;
		Addr <=  "0101000101010";
		Trees_din <= x"ff792a19";
		wait for Clk_period;
		Addr <=  "0101000101011";
		Trees_din <= x"fff12a19";
		wait for Clk_period;
		Addr <=  "0101000101100";
		Trees_din <= x"d8000304";
		wait for Clk_period;
		Addr <=  "0101000101101";
		Trees_din <= x"ffc32a19";
		wait for Clk_period;
		Addr <=  "0101000101110";
		Trees_din <= x"76ffff04";
		wait for Clk_period;
		Addr <=  "0101000101111";
		Trees_din <= x"009d2a19";
		wait for Clk_period;
		Addr <=  "0101000110000";
		Trees_din <= x"001f2a19";
		wait for Clk_period;
		Addr <=  "0101000110001";
		Trees_din <= x"19ff8110";
		wait for Clk_period;
		Addr <=  "0101000110010";
		Trees_din <= x"57ff3608";
		wait for Clk_period;
		Addr <=  "0101000110011";
		Trees_din <= x"e7ffdf04";
		wait for Clk_period;
		Addr <=  "0101000110100";
		Trees_din <= x"ff922a19";
		wait for Clk_period;
		Addr <=  "0101000110101";
		Trees_din <= x"fff82a19";
		wait for Clk_period;
		Addr <=  "0101000110110";
		Trees_din <= x"d2feca04";
		wait for Clk_period;
		Addr <=  "0101000110111";
		Trees_din <= x"004c2a19";
		wait for Clk_period;
		Addr <=  "0101000111000";
		Trees_din <= x"ffad2a19";
		wait for Clk_period;
		Addr <=  "0101000111001";
		Trees_din <= x"7cffa408";
		wait for Clk_period;
		Addr <=  "0101000111010";
		Trees_din <= x"77fe9404";
		wait for Clk_period;
		Addr <=  "0101000111011";
		Trees_din <= x"00452a19";
		wait for Clk_period;
		Addr <=  "0101000111100";
		Trees_din <= x"ff972a19";
		wait for Clk_period;
		Addr <=  "0101000111101";
		Trees_din <= x"66ffea04";
		wait for Clk_period;
		Addr <=  "0101000111110";
		Trees_din <= x"008c2a19";
		wait for Clk_period;
		Addr <=  "0101000111111";
		Trees_din <= x"fffb2a19";
		wait for Clk_period;
		Addr <=  "0101001000000";
		Trees_din <= x"7dff771c";
		wait for Clk_period;
		Addr <=  "0101001000001";
		Trees_din <= x"b6ff710c";
		wait for Clk_period;
		Addr <=  "0101001000010";
		Trees_din <= x"f3003308";
		wait for Clk_period;
		Addr <=  "0101001000011";
		Trees_din <= x"82001e04";
		wait for Clk_period;
		Addr <=  "0101001000100";
		Trees_din <= x"00482a19";
		wait for Clk_period;
		Addr <=  "0101001000101";
		Trees_din <= x"ffbc2a19";
		wait for Clk_period;
		Addr <=  "0101001000110";
		Trees_din <= x"ff6c2a19";
		wait for Clk_period;
		Addr <=  "0101001000111";
		Trees_din <= x"2cff8108";
		wait for Clk_period;
		Addr <=  "0101001001000";
		Trees_din <= x"9eff4504";
		wait for Clk_period;
		Addr <=  "0101001001001";
		Trees_din <= x"001f2a19";
		wait for Clk_period;
		Addr <=  "0101001001010";
		Trees_din <= x"ff6f2a19";
		wait for Clk_period;
		Addr <=  "0101001001011";
		Trees_din <= x"72ffe204";
		wait for Clk_period;
		Addr <=  "0101001001100";
		Trees_din <= x"00732a19";
		wait for Clk_period;
		Addr <=  "0101001001101";
		Trees_din <= x"ffe02a19";
		wait for Clk_period;
		Addr <=  "0101001001110";
		Trees_din <= x"9dffc910";
		wait for Clk_period;
		Addr <=  "0101001001111";
		Trees_din <= x"da000b08";
		wait for Clk_period;
		Addr <=  "0101001010000";
		Trees_din <= x"d600af04";
		wait for Clk_period;
		Addr <=  "0101001010001";
		Trees_din <= x"001e2a19";
		wait for Clk_period;
		Addr <=  "0101001010010";
		Trees_din <= x"ffb62a19";
		wait for Clk_period;
		Addr <=  "0101001010011";
		Trees_din <= x"edff9d04";
		wait for Clk_period;
		Addr <=  "0101001010100";
		Trees_din <= x"001c2a19";
		wait for Clk_period;
		Addr <=  "0101001010101";
		Trees_din <= x"ffc42a19";
		wait for Clk_period;
		Addr <=  "0101001010110";
		Trees_din <= x"53ffa708";
		wait for Clk_period;
		Addr <=  "0101001010111";
		Trees_din <= x"bfffc804";
		wait for Clk_period;
		Addr <=  "0101001011000";
		Trees_din <= x"ffe32a19";
		wait for Clk_period;
		Addr <=  "0101001011001";
		Trees_din <= x"00422a19";
		wait for Clk_period;
		Addr <=  "0101001011010";
		Trees_din <= x"03ff4a04";
		wait for Clk_period;
		Addr <=  "0101001011011";
		Trees_din <= x"002e2a19";
		wait for Clk_period;
		Addr <=  "0101001011100";
		Trees_din <= x"ffa02a19";
		wait for Clk_period;
		Addr <=  "0101001011101";
		Trees_din <= x"21ff6820";
		wait for Clk_period;
		Addr <=  "0101001011110";
		Trees_din <= x"edff1808";
		wait for Clk_period;
		Addr <=  "0101001011111";
		Trees_din <= x"c3003004";
		wait for Clk_period;
		Addr <=  "0101001100000";
		Trees_din <= x"00812a19";
		wait for Clk_period;
		Addr <=  "0101001100001";
		Trees_din <= x"ffdb2a19";
		wait for Clk_period;
		Addr <=  "0101001100010";
		Trees_din <= x"d7009410";
		wait for Clk_period;
		Addr <=  "0101001100011";
		Trees_din <= x"a2ff9808";
		wait for Clk_period;
		Addr <=  "0101001100100";
		Trees_din <= x"f1ffab04";
		wait for Clk_period;
		Addr <=  "0101001100101";
		Trees_din <= x"ff762a19";
		wait for Clk_period;
		Addr <=  "0101001100110";
		Trees_din <= x"00452a19";
		wait for Clk_period;
		Addr <=  "0101001100111";
		Trees_din <= x"70fe8f04";
		wait for Clk_period;
		Addr <=  "0101001101000";
		Trees_din <= x"ffb42a19";
		wait for Clk_period;
		Addr <=  "0101001101001";
		Trees_din <= x"00652a19";
		wait for Clk_period;
		Addr <=  "0101001101010";
		Trees_din <= x"0d001104";
		wait for Clk_period;
		Addr <=  "0101001101011";
		Trees_din <= x"ff5c2a19";
		wait for Clk_period;
		Addr <=  "0101001101100";
		Trees_din <= x"00022a19";
		wait for Clk_period;
		Addr <=  "0101001101101";
		Trees_din <= x"49ffa61c";
		wait for Clk_period;
		Addr <=  "0101001101110";
		Trees_din <= x"e0fed70c";
		wait for Clk_period;
		Addr <=  "0101001101111";
		Trees_din <= x"46feab04";
		wait for Clk_period;
		Addr <=  "0101001110000";
		Trees_din <= x"00332a19";
		wait for Clk_period;
		Addr <=  "0101001110001";
		Trees_din <= x"67ffc804";
		wait for Clk_period;
		Addr <=  "0101001110010";
		Trees_din <= x"ff742a19";
		wait for Clk_period;
		Addr <=  "0101001110011";
		Trees_din <= x"000a2a19";
		wait for Clk_period;
		Addr <=  "0101001110100";
		Trees_din <= x"baffc708";
		wait for Clk_period;
		Addr <=  "0101001110101";
		Trees_din <= x"c6ff5504";
		wait for Clk_period;
		Addr <=  "0101001110110";
		Trees_din <= x"ff8a2a19";
		wait for Clk_period;
		Addr <=  "0101001110111";
		Trees_din <= x"002d2a19";
		wait for Clk_period;
		Addr <=  "0101001111000";
		Trees_din <= x"d3ff6904";
		wait for Clk_period;
		Addr <=  "0101001111001";
		Trees_din <= x"007c2a19";
		wait for Clk_period;
		Addr <=  "0101001111010";
		Trees_din <= x"ffd02a19";
		wait for Clk_period;
		Addr <=  "0101001111011";
		Trees_din <= x"da00a410";
		wait for Clk_period;
		Addr <=  "0101001111100";
		Trees_din <= x"4dfdb508";
		wait for Clk_period;
		Addr <=  "0101001111101";
		Trees_din <= x"4cfe6c04";
		wait for Clk_period;
		Addr <=  "0101001111110";
		Trees_din <= x"00312a19";
		wait for Clk_period;
		Addr <=  "0101001111111";
		Trees_din <= x"ff6e2a19";
		wait for Clk_period;
		Addr <=  "0101010000000";
		Trees_din <= x"e1007d04";
		wait for Clk_period;
		Addr <=  "0101010000001";
		Trees_din <= x"00452a19";
		wait for Clk_period;
		Addr <=  "0101010000010";
		Trees_din <= x"ff9c2a19";
		wait for Clk_period;
		Addr <=  "0101010000011";
		Trees_din <= x"40ffd104";
		wait for Clk_period;
		Addr <=  "0101010000100";
		Trees_din <= x"00292a19";
		wait for Clk_period;
		Addr <=  "0101010000101";
		Trees_din <= x"ff7f2a19";
		wait for Clk_period;
		Addr <=  "0101010000110";
		Trees_din <= x"1efef228";
		wait for Clk_period;
		Addr <=  "0101010000111";
		Trees_din <= x"2400091c";
		wait for Clk_period;
		Addr <=  "0101010001000";
		Trees_din <= x"84ff420c";
		wait for Clk_period;
		Addr <=  "0101010001001";
		Trees_din <= x"0800ac08";
		wait for Clk_period;
		Addr <=  "0101010001010";
		Trees_din <= x"56ff8604";
		wait for Clk_period;
		Addr <=  "0101010001011";
		Trees_din <= x"00052b65";
		wait for Clk_period;
		Addr <=  "0101010001100";
		Trees_din <= x"006e2b65";
		wait for Clk_period;
		Addr <=  "0101010001101";
		Trees_din <= x"ffbe2b65";
		wait for Clk_period;
		Addr <=  "0101010001110";
		Trees_din <= x"93fea404";
		wait for Clk_period;
		Addr <=  "0101010001111";
		Trees_din <= x"003b2b65";
		wait for Clk_period;
		Addr <=  "0101010010000";
		Trees_din <= x"cfffb904";
		wait for Clk_period;
		Addr <=  "0101010010001";
		Trees_din <= x"00112b65";
		wait for Clk_period;
		Addr <=  "0101010010010";
		Trees_din <= x"3d005504";
		wait for Clk_period;
		Addr <=  "0101010010011";
		Trees_din <= x"ff652b65";
		wait for Clk_period;
		Addr <=  "0101010010100";
		Trees_din <= x"ffe72b65";
		wait for Clk_period;
		Addr <=  "0101010010101";
		Trees_din <= x"60ffa708";
		wait for Clk_period;
		Addr <=  "0101010010110";
		Trees_din <= x"40002504";
		wait for Clk_period;
		Addr <=  "0101010010111";
		Trees_din <= x"00802b65";
		wait for Clk_period;
		Addr <=  "0101010011000";
		Trees_din <= x"ffe62b65";
		wait for Clk_period;
		Addr <=  "0101010011001";
		Trees_din <= x"ffc12b65";
		wait for Clk_period;
		Addr <=  "0101010011010";
		Trees_din <= x"09ffe240";
		wait for Clk_period;
		Addr <=  "0101010011011";
		Trees_din <= x"1fff7720";
		wait for Clk_period;
		Addr <=  "0101010011100";
		Trees_din <= x"dc003c10";
		wait for Clk_period;
		Addr <=  "0101010011101";
		Trees_din <= x"6bfe3408";
		wait for Clk_period;
		Addr <=  "0101010011110";
		Trees_din <= x"3d000004";
		wait for Clk_period;
		Addr <=  "0101010011111";
		Trees_din <= x"00312b65";
		wait for Clk_period;
		Addr <=  "0101010100000";
		Trees_din <= x"ff8f2b65";
		wait for Clk_period;
		Addr <=  "0101010100001";
		Trees_din <= x"8fff7404";
		wait for Clk_period;
		Addr <=  "0101010100010";
		Trees_din <= x"00422b65";
		wait for Clk_period;
		Addr <=  "0101010100011";
		Trees_din <= x"ffdf2b65";
		wait for Clk_period;
		Addr <=  "0101010100100";
		Trees_din <= x"59ffc408";
		wait for Clk_period;
		Addr <=  "0101010100101";
		Trees_din <= x"e4ff2504";
		wait for Clk_period;
		Addr <=  "0101010100110";
		Trees_din <= x"ff932b65";
		wait for Clk_period;
		Addr <=  "0101010100111";
		Trees_din <= x"00392b65";
		wait for Clk_period;
		Addr <=  "0101010101000";
		Trees_din <= x"c7fead04";
		wait for Clk_period;
		Addr <=  "0101010101001";
		Trees_din <= x"ffad2b65";
		wait for Clk_period;
		Addr <=  "0101010101010";
		Trees_din <= x"00782b65";
		wait for Clk_period;
		Addr <=  "0101010101011";
		Trees_din <= x"71000d10";
		wait for Clk_period;
		Addr <=  "0101010101100";
		Trees_din <= x"45ff0808";
		wait for Clk_period;
		Addr <=  "0101010101101";
		Trees_din <= x"d6004c04";
		wait for Clk_period;
		Addr <=  "0101010101110";
		Trees_din <= x"00022b65";
		wait for Clk_period;
		Addr <=  "0101010101111";
		Trees_din <= x"ffc32b65";
		wait for Clk_period;
		Addr <=  "0101010110000";
		Trees_din <= x"2bff3d04";
		wait for Clk_period;
		Addr <=  "0101010110001";
		Trees_din <= x"ffbe2b65";
		wait for Clk_period;
		Addr <=  "0101010110010";
		Trees_din <= x"00272b65";
		wait for Clk_period;
		Addr <=  "0101010110011";
		Trees_din <= x"be005a08";
		wait for Clk_period;
		Addr <=  "0101010110100";
		Trees_din <= x"65ffcc04";
		wait for Clk_period;
		Addr <=  "0101010110101";
		Trees_din <= x"ff7b2b65";
		wait for Clk_period;
		Addr <=  "0101010110110";
		Trees_din <= x"00222b65";
		wait for Clk_period;
		Addr <=  "0101010110111";
		Trees_din <= x"2eff9a04";
		wait for Clk_period;
		Addr <=  "0101010111000";
		Trees_din <= x"00642b65";
		wait for Clk_period;
		Addr <=  "0101010111001";
		Trees_din <= x"fffb2b65";
		wait for Clk_period;
		Addr <=  "0101010111010";
		Trees_din <= x"5bffa120";
		wait for Clk_period;
		Addr <=  "0101010111011";
		Trees_din <= x"d2fee810";
		wait for Clk_period;
		Addr <=  "0101010111100";
		Trees_din <= x"25ffd908";
		wait for Clk_period;
		Addr <=  "0101010111101";
		Trees_din <= x"d8005104";
		wait for Clk_period;
		Addr <=  "0101010111110";
		Trees_din <= x"005d2b65";
		wait for Clk_period;
		Addr <=  "0101010111111";
		Trees_din <= x"ffc62b65";
		wait for Clk_period;
		Addr <=  "0101011000000";
		Trees_din <= x"35fe7604";
		wait for Clk_period;
		Addr <=  "0101011000001";
		Trees_din <= x"00202b65";
		wait for Clk_period;
		Addr <=  "0101011000010";
		Trees_din <= x"ffca2b65";
		wait for Clk_period;
		Addr <=  "0101011000011";
		Trees_din <= x"77fe9e08";
		wait for Clk_period;
		Addr <=  "0101011000100";
		Trees_din <= x"aefef504";
		wait for Clk_period;
		Addr <=  "0101011000101";
		Trees_din <= x"ffab2b65";
		wait for Clk_period;
		Addr <=  "0101011000110";
		Trees_din <= x"00622b65";
		wait for Clk_period;
		Addr <=  "0101011000111";
		Trees_din <= x"98fe1604";
		wait for Clk_period;
		Addr <=  "0101011001000";
		Trees_din <= x"00612b65";
		wait for Clk_period;
		Addr <=  "0101011001001";
		Trees_din <= x"ff9c2b65";
		wait for Clk_period;
		Addr <=  "0101011001010";
		Trees_din <= x"76ffc210";
		wait for Clk_period;
		Addr <=  "0101011001011";
		Trees_din <= x"4bff2e08";
		wait for Clk_period;
		Addr <=  "0101011001100";
		Trees_din <= x"96feed04";
		wait for Clk_period;
		Addr <=  "0101011001101";
		Trees_din <= x"fff72b65";
		wait for Clk_period;
		Addr <=  "0101011001110";
		Trees_din <= x"00862b65";
		wait for Clk_period;
		Addr <=  "0101011001111";
		Trees_din <= x"dbffdc04";
		wait for Clk_period;
		Addr <=  "0101011010000";
		Trees_din <= x"ff8e2b65";
		wait for Clk_period;
		Addr <=  "0101011010001";
		Trees_din <= x"00312b65";
		wait for Clk_period;
		Addr <=  "0101011010010";
		Trees_din <= x"eaffb208";
		wait for Clk_period;
		Addr <=  "0101011010011";
		Trees_din <= x"1cff2d04";
		wait for Clk_period;
		Addr <=  "0101011010100";
		Trees_din <= x"003f2b65";
		wait for Clk_period;
		Addr <=  "0101011010101";
		Trees_din <= x"ff922b65";
		wait for Clk_period;
		Addr <=  "0101011010110";
		Trees_din <= x"a4ff9d04";
		wait for Clk_period;
		Addr <=  "0101011010111";
		Trees_din <= x"001f2b65";
		wait for Clk_period;
		Addr <=  "0101011011000";
		Trees_din <= x"00802b65";
		wait for Clk_period;
		Addr <=  "0101011011001";
		Trees_din <= x"3100b660";
		wait for Clk_period;
		Addr <=  "0101011011010";
		Trees_din <= x"43ffa738";
		wait for Clk_period;
		Addr <=  "0101011011011";
		Trees_din <= x"a1000e20";
		wait for Clk_period;
		Addr <=  "0101011011100";
		Trees_din <= x"b2ffa410";
		wait for Clk_period;
		Addr <=  "0101011011101";
		Trees_din <= x"ecffff08";
		wait for Clk_period;
		Addr <=  "0101011011110";
		Trees_din <= x"a5ff6c04";
		wait for Clk_period;
		Addr <=  "0101011011111";
		Trees_din <= x"00092c61";
		wait for Clk_period;
		Addr <=  "0101011100000";
		Trees_din <= x"ff9d2c61";
		wait for Clk_period;
		Addr <=  "0101011100001";
		Trees_din <= x"e0ff9504";
		wait for Clk_period;
		Addr <=  "0101011100010";
		Trees_din <= x"ff9b2c61";
		wait for Clk_period;
		Addr <=  "0101011100011";
		Trees_din <= x"00132c61";
		wait for Clk_period;
		Addr <=  "0101011100100";
		Trees_din <= x"58ff1108";
		wait for Clk_period;
		Addr <=  "0101011100101";
		Trees_din <= x"02feb304";
		wait for Clk_period;
		Addr <=  "0101011100110";
		Trees_din <= x"000a2c61";
		wait for Clk_period;
		Addr <=  "0101011100111";
		Trees_din <= x"ffdd2c61";
		wait for Clk_period;
		Addr <=  "0101011101000";
		Trees_din <= x"5c003204";
		wait for Clk_period;
		Addr <=  "0101011101001";
		Trees_din <= x"00302c61";
		wait for Clk_period;
		Addr <=  "0101011101010";
		Trees_din <= x"fff12c61";
		wait for Clk_period;
		Addr <=  "0101011101011";
		Trees_din <= x"2bffab10";
		wait for Clk_period;
		Addr <=  "0101011101100";
		Trees_din <= x"a5ff4308";
		wait for Clk_period;
		Addr <=  "0101011101101";
		Trees_din <= x"1bffa804";
		wait for Clk_period;
		Addr <=  "0101011101110";
		Trees_din <= x"00752c61";
		wait for Clk_period;
		Addr <=  "0101011101111";
		Trees_din <= x"fff02c61";
		wait for Clk_period;
		Addr <=  "0101011110000";
		Trees_din <= x"15ff3e04";
		wait for Clk_period;
		Addr <=  "0101011110001";
		Trees_din <= x"fff62c61";
		wait for Clk_period;
		Addr <=  "0101011110010";
		Trees_din <= x"ff8a2c61";
		wait for Clk_period;
		Addr <=  "0101011110011";
		Trees_din <= x"eaffe204";
		wait for Clk_period;
		Addr <=  "0101011110100";
		Trees_din <= x"00942c61";
		wait for Clk_period;
		Addr <=  "0101011110101";
		Trees_din <= x"00202c61";
		wait for Clk_period;
		Addr <=  "0101011110110";
		Trees_din <= x"06fed308";
		wait for Clk_period;
		Addr <=  "0101011110111";
		Trees_din <= x"90ff1004";
		wait for Clk_period;
		Addr <=  "0101011111000";
		Trees_din <= x"00212c61";
		wait for Clk_period;
		Addr <=  "0101011111001";
		Trees_din <= x"ff7d2c61";
		wait for Clk_period;
		Addr <=  "0101011111010";
		Trees_din <= x"44ffe110";
		wait for Clk_period;
		Addr <=  "0101011111011";
		Trees_din <= x"b3ff7308";
		wait for Clk_period;
		Addr <=  "0101011111100";
		Trees_din <= x"36fe9704";
		wait for Clk_period;
		Addr <=  "0101011111101";
		Trees_din <= x"ffbc2c61";
		wait for Clk_period;
		Addr <=  "0101011111110";
		Trees_din <= x"00502c61";
		wait for Clk_period;
		Addr <=  "0101011111111";
		Trees_din <= x"ecffef04";
		wait for Clk_period;
		Addr <=  "0101100000000";
		Trees_din <= x"ff872c61";
		wait for Clk_period;
		Addr <=  "0101100000001";
		Trees_din <= x"004f2c61";
		wait for Clk_period;
		Addr <=  "0101100000010";
		Trees_din <= x"ddfede08";
		wait for Clk_period;
		Addr <=  "0101100000011";
		Trees_din <= x"1dfe9604";
		wait for Clk_period;
		Addr <=  "0101100000100";
		Trees_din <= x"00472c61";
		wait for Clk_period;
		Addr <=  "0101100000101";
		Trees_din <= x"ff9f2c61";
		wait for Clk_period;
		Addr <=  "0101100000110";
		Trees_din <= x"49ffa904";
		wait for Clk_period;
		Addr <=  "0101100000111";
		Trees_din <= x"ffd52c61";
		wait for Clk_period;
		Addr <=  "0101100001000";
		Trees_din <= x"002a2c61";
		wait for Clk_period;
		Addr <=  "0101100001001";
		Trees_din <= x"4bfe3004";
		wait for Clk_period;
		Addr <=  "0101100001010";
		Trees_din <= x"00532c61";
		wait for Clk_period;
		Addr <=  "0101100001011";
		Trees_din <= x"cffff80c";
		wait for Clk_period;
		Addr <=  "0101100001100";
		Trees_din <= x"c9ff9804";
		wait for Clk_period;
		Addr <=  "0101100001101";
		Trees_din <= x"ffa62c61";
		wait for Clk_period;
		Addr <=  "0101100001110";
		Trees_din <= x"33ff2b04";
		wait for Clk_period;
		Addr <=  "0101100001111";
		Trees_din <= x"ffcb2c61";
		wait for Clk_period;
		Addr <=  "0101100010000";
		Trees_din <= x"00742c61";
		wait for Clk_period;
		Addr <=  "0101100010001";
		Trees_din <= x"7eff2a0c";
		wait for Clk_period;
		Addr <=  "0101100010010";
		Trees_din <= x"1e000f08";
		wait for Clk_period;
		Addr <=  "0101100010011";
		Trees_din <= x"6effaf04";
		wait for Clk_period;
		Addr <=  "0101100010100";
		Trees_din <= x"00062c61";
		wait for Clk_period;
		Addr <=  "0101100010101";
		Trees_din <= x"ff642c61";
		wait for Clk_period;
		Addr <=  "0101100010110";
		Trees_din <= x"001a2c61";
		wait for Clk_period;
		Addr <=  "0101100010111";
		Trees_din <= x"000f2c61";
		wait for Clk_period;
		Addr <=  "0101100011000";
		Trees_din <= x"f5007e74";
		wait for Clk_period;
		Addr <=  "0101100011001";
		Trees_din <= x"8fff343c";
		wait for Clk_period;
		Addr <=  "0101100011010";
		Trees_din <= x"b6fe8d1c";
		wait for Clk_period;
		Addr <=  "0101100011011";
		Trees_din <= x"a9ff630c";
		wait for Clk_period;
		Addr <=  "0101100011100";
		Trees_din <= x"2bffbd04";
		wait for Clk_period;
		Addr <=  "0101100011101";
		Trees_din <= x"007f2d85";
		wait for Clk_period;
		Addr <=  "0101100011110";
		Trees_din <= x"77fe7004";
		wait for Clk_period;
		Addr <=  "0101100011111";
		Trees_din <= x"ff9b2d85";
		wait for Clk_period;
		Addr <=  "0101100100000";
		Trees_din <= x"ffff2d85";
		wait for Clk_period;
		Addr <=  "0101100100001";
		Trees_din <= x"b1ff1808";
		wait for Clk_period;
		Addr <=  "0101100100010";
		Trees_din <= x"8cff5704";
		wait for Clk_period;
		Addr <=  "0101100100011";
		Trees_din <= x"fff82d85";
		wait for Clk_period;
		Addr <=  "0101100100100";
		Trees_din <= x"ff4e2d85";
		wait for Clk_period;
		Addr <=  "0101100100101";
		Trees_din <= x"7affd504";
		wait for Clk_period;
		Addr <=  "0101100100110";
		Trees_din <= x"00352d85";
		wait for Clk_period;
		Addr <=  "0101100100111";
		Trees_din <= x"ff872d85";
		wait for Clk_period;
		Addr <=  "0101100101000";
		Trees_din <= x"a8ff2810";
		wait for Clk_period;
		Addr <=  "0101100101001";
		Trees_din <= x"fcff3e08";
		wait for Clk_period;
		Addr <=  "0101100101010";
		Trees_din <= x"64ffef04";
		wait for Clk_period;
		Addr <=  "0101100101011";
		Trees_din <= x"00152d85";
		wait for Clk_period;
		Addr <=  "0101100101100";
		Trees_din <= x"ff8a2d85";
		wait for Clk_period;
		Addr <=  "0101100101101";
		Trees_din <= x"20ffeb04";
		wait for Clk_period;
		Addr <=  "0101100101110";
		Trees_din <= x"ffe92d85";
		wait for Clk_period;
		Addr <=  "0101100101111";
		Trees_din <= x"ff882d85";
		wait for Clk_period;
		Addr <=  "0101100110000";
		Trees_din <= x"91ff7508";
		wait for Clk_period;
		Addr <=  "0101100110001";
		Trees_din <= x"24ff9c04";
		wait for Clk_period;
		Addr <=  "0101100110010";
		Trees_din <= x"ffd82d85";
		wait for Clk_period;
		Addr <=  "0101100110011";
		Trees_din <= x"00102d85";
		wait for Clk_period;
		Addr <=  "0101100110100";
		Trees_din <= x"3dffaa04";
		wait for Clk_period;
		Addr <=  "0101100110101";
		Trees_din <= x"fff52d85";
		wait for Clk_period;
		Addr <=  "0101100110110";
		Trees_din <= x"002f2d85";
		wait for Clk_period;
		Addr <=  "0101100110111";
		Trees_din <= x"01fec31c";
		wait for Clk_period;
		Addr <=  "0101100111000";
		Trees_din <= x"e1ff680c";
		wait for Clk_period;
		Addr <=  "0101100111001";
		Trees_din <= x"a0fe0404";
		wait for Clk_period;
		Addr <=  "0101100111010";
		Trees_din <= x"ff802d85";
		wait for Clk_period;
		Addr <=  "0101100111011";
		Trees_din <= x"59ff9904";
		wait for Clk_period;
		Addr <=  "0101100111100";
		Trees_din <= x"ffd92d85";
		wait for Clk_period;
		Addr <=  "0101100111101";
		Trees_din <= x"005a2d85";
		wait for Clk_period;
		Addr <=  "0101100111110";
		Trees_din <= x"b7ff5208";
		wait for Clk_period;
		Addr <=  "0101100111111";
		Trees_din <= x"12ffdc04";
		wait for Clk_period;
		Addr <=  "0101101000000";
		Trees_din <= x"00542d85";
		wait for Clk_period;
		Addr <=  "0101101000001";
		Trees_din <= x"ffb52d85";
		wait for Clk_period;
		Addr <=  "0101101000010";
		Trees_din <= x"c9ff3304";
		wait for Clk_period;
		Addr <=  "0101101000011";
		Trees_din <= x"00532d85";
		wait for Clk_period;
		Addr <=  "0101101000100";
		Trees_din <= x"ffa72d85";
		wait for Clk_period;
		Addr <=  "0101101000101";
		Trees_din <= x"97ff7b10";
		wait for Clk_period;
		Addr <=  "0101101000110";
		Trees_din <= x"53ff6208";
		wait for Clk_period;
		Addr <=  "0101101000111";
		Trees_din <= x"60ff2004";
		wait for Clk_period;
		Addr <=  "0101101001000";
		Trees_din <= x"ffdb2d85";
		wait for Clk_period;
		Addr <=  "0101101001001";
		Trees_din <= x"00652d85";
		wait for Clk_period;
		Addr <=  "0101101001010";
		Trees_din <= x"6d001b04";
		wait for Clk_period;
		Addr <=  "0101101001011";
		Trees_din <= x"00282d85";
		wait for Clk_period;
		Addr <=  "0101101001100";
		Trees_din <= x"ffc02d85";
		wait for Clk_period;
		Addr <=  "0101101001101";
		Trees_din <= x"aaff0e04";
		wait for Clk_period;
		Addr <=  "0101101001110";
		Trees_din <= x"00652d85";
		wait for Clk_period;
		Addr <=  "0101101001111";
		Trees_din <= x"32fe9a04";
		wait for Clk_period;
		Addr <=  "0101101010000";
		Trees_din <= x"004a2d85";
		wait for Clk_period;
		Addr <=  "0101101010001";
		Trees_din <= x"ffaa2d85";
		wait for Clk_period;
		Addr <=  "0101101010010";
		Trees_din <= x"2dff4318";
		wait for Clk_period;
		Addr <=  "0101101010011";
		Trees_din <= x"bf000f10";
		wait for Clk_period;
		Addr <=  "0101101010100";
		Trees_din <= x"ee00c40c";
		wait for Clk_period;
		Addr <=  "0101101010101";
		Trees_din <= x"70ff8e08";
		wait for Clk_period;
		Addr <=  "0101101010110";
		Trees_din <= x"cd000104";
		wait for Clk_period;
		Addr <=  "0101101010111";
		Trees_din <= x"00902d85";
		wait for Clk_period;
		Addr <=  "0101101011000";
		Trees_din <= x"001c2d85";
		wait for Clk_period;
		Addr <=  "0101101011001";
		Trees_din <= x"ffe22d85";
		wait for Clk_period;
		Addr <=  "0101101011010";
		Trees_din <= x"ffd02d85";
		wait for Clk_period;
		Addr <=  "0101101011011";
		Trees_din <= x"cdffb004";
		wait for Clk_period;
		Addr <=  "0101101011100";
		Trees_din <= x"ff932d85";
		wait for Clk_period;
		Addr <=  "0101101011101";
		Trees_din <= x"00032d85";
		wait for Clk_period;
		Addr <=  "0101101011110";
		Trees_din <= x"04001104";
		wait for Clk_period;
		Addr <=  "0101101011111";
		Trees_din <= x"00112d85";
		wait for Clk_period;
		Addr <=  "0101101100000";
		Trees_din <= x"ffa12d85";
		wait for Clk_period;
		Addr <=  "0101101100001";
		Trees_din <= x"7c01097c";
		wait for Clk_period;
		Addr <=  "0101101100010";
		Trees_din <= x"6d003c3c";
		wait for Clk_period;
		Addr <=  "0101101100011";
		Trees_din <= x"a4ff081c";
		wait for Clk_period;
		Addr <=  "0101101100100";
		Trees_din <= x"9afff210";
		wait for Clk_period;
		Addr <=  "0101101100101";
		Trees_din <= x"47ffab08";
		wait for Clk_period;
		Addr <=  "0101101100110";
		Trees_din <= x"c5ff0604";
		wait for Clk_period;
		Addr <=  "0101101100111";
		Trees_din <= x"ffe32e89";
		wait for Clk_period;
		Addr <=  "0101101101000";
		Trees_din <= x"00732e89";
		wait for Clk_period;
		Addr <=  "0101101101001";
		Trees_din <= x"ceffb004";
		wait for Clk_period;
		Addr <=  "0101101101010";
		Trees_din <= x"ff902e89";
		wait for Clk_period;
		Addr <=  "0101101101011";
		Trees_din <= x"00232e89";
		wait for Clk_period;
		Addr <=  "0101101101100";
		Trees_din <= x"c8001c08";
		wait for Clk_period;
		Addr <=  "0101101101101";
		Trees_din <= x"e3ff0004";
		wait for Clk_period;
		Addr <=  "0101101101110";
		Trees_din <= x"ff622e89";
		wait for Clk_period;
		Addr <=  "0101101101111";
		Trees_din <= x"00132e89";
		wait for Clk_period;
		Addr <=  "0101101110000";
		Trees_din <= x"004b2e89";
		wait for Clk_period;
		Addr <=  "0101101110001";
		Trees_din <= x"21000110";
		wait for Clk_period;
		Addr <=  "0101101110010";
		Trees_din <= x"9bfebf08";
		wait for Clk_period;
		Addr <=  "0101101110011";
		Trees_din <= x"fdff5204";
		wait for Clk_period;
		Addr <=  "0101101110100";
		Trees_din <= x"00122e89";
		wait for Clk_period;
		Addr <=  "0101101110101";
		Trees_din <= x"ffb22e89";
		wait for Clk_period;
		Addr <=  "0101101110110";
		Trees_din <= x"50ff6f04";
		wait for Clk_period;
		Addr <=  "0101101110111";
		Trees_din <= x"fff52e89";
		wait for Clk_period;
		Addr <=  "0101101111000";
		Trees_din <= x"001b2e89";
		wait for Clk_period;
		Addr <=  "0101101111001";
		Trees_din <= x"6e009d08";
		wait for Clk_period;
		Addr <=  "0101101111010";
		Trees_din <= x"72006b04";
		wait for Clk_period;
		Addr <=  "0101101111011";
		Trees_din <= x"004a2e89";
		wait for Clk_period;
		Addr <=  "0101101111100";
		Trees_din <= x"fff22e89";
		wait for Clk_period;
		Addr <=  "0101101111101";
		Trees_din <= x"76ffd704";
		wait for Clk_period;
		Addr <=  "0101101111110";
		Trees_din <= x"00172e89";
		wait for Clk_period;
		Addr <=  "0101101111111";
		Trees_din <= x"ff822e89";
		wait for Clk_period;
		Addr <=  "0101110000000";
		Trees_din <= x"ee003b20";
		wait for Clk_period;
		Addr <=  "0101110000001";
		Trees_din <= x"45ff1e10";
		wait for Clk_period;
		Addr <=  "0101110000010";
		Trees_din <= x"f2038708";
		wait for Clk_period;
		Addr <=  "0101110000011";
		Trees_din <= x"59000904";
		wait for Clk_period;
		Addr <=  "0101110000100";
		Trees_din <= x"ffb32e89";
		wait for Clk_period;
		Addr <=  "0101110000101";
		Trees_din <= x"fff92e89";
		wait for Clk_period;
		Addr <=  "0101110000110";
		Trees_din <= x"ebfea104";
		wait for Clk_period;
		Addr <=  "0101110000111";
		Trees_din <= x"ffd62e89";
		wait for Clk_period;
		Addr <=  "0101110001000";
		Trees_din <= x"00712e89";
		wait for Clk_period;
		Addr <=  "0101110001001";
		Trees_din <= x"0dff9608";
		wait for Clk_period;
		Addr <=  "0101110001010";
		Trees_din <= x"3d000e04";
		wait for Clk_period;
		Addr <=  "0101110001011";
		Trees_din <= x"00132e89";
		wait for Clk_period;
		Addr <=  "0101110001100";
		Trees_din <= x"ffa82e89";
		wait for Clk_period;
		Addr <=  "0101110001101";
		Trees_din <= x"0b004904";
		wait for Clk_period;
		Addr <=  "0101110001110";
		Trees_din <= x"00612e89";
		wait for Clk_period;
		Addr <=  "0101110001111";
		Trees_din <= x"ffc42e89";
		wait for Clk_period;
		Addr <=  "0101110010000";
		Trees_din <= x"20ff3710";
		wait for Clk_period;
		Addr <=  "0101110010001";
		Trees_din <= x"23ff0d08";
		wait for Clk_period;
		Addr <=  "0101110010010";
		Trees_din <= x"23fef404";
		wait for Clk_period;
		Addr <=  "0101110010011";
		Trees_din <= x"00442e89";
		wait for Clk_period;
		Addr <=  "0101110010100";
		Trees_din <= x"ff992e89";
		wait for Clk_period;
		Addr <=  "0101110010101";
		Trees_din <= x"81ff7104";
		wait for Clk_period;
		Addr <=  "0101110010110";
		Trees_din <= x"001a2e89";
		wait for Clk_period;
		Addr <=  "0101110010111";
		Trees_din <= x"00892e89";
		wait for Clk_period;
		Addr <=  "0101110011000";
		Trees_din <= x"01fe6408";
		wait for Clk_period;
		Addr <=  "0101110011001";
		Trees_din <= x"32fef504";
		wait for Clk_period;
		Addr <=  "0101110011010";
		Trees_din <= x"ff7f2e89";
		wait for Clk_period;
		Addr <=  "0101110011011";
		Trees_din <= x"00312e89";
		wait for Clk_period;
		Addr <=  "0101110011100";
		Trees_din <= x"c7ff0204";
		wait for Clk_period;
		Addr <=  "0101110011101";
		Trees_din <= x"fff52e89";
		wait for Clk_period;
		Addr <=  "0101110011110";
		Trees_din <= x"00522e89";
		wait for Clk_period;
		Addr <=  "0101110011111";
		Trees_din <= x"0cfe0304";
		wait for Clk_period;
		Addr <=  "0101110100000";
		Trees_din <= x"ffcc2e89";
		wait for Clk_period;
		Addr <=  "0101110100001";
		Trees_din <= x"00902e89";
		wait for Clk_period;
		Addr <=  "0101110100010";
		Trees_din <= x"7d00456c";
		wait for Clk_period;
		Addr <=  "0101110100011";
		Trees_din <= x"31feff30";
		wait for Clk_period;
		Addr <=  "0101110100100";
		Trees_din <= x"20ff6c18";
		wait for Clk_period;
		Addr <=  "0101110100101";
		Trees_din <= x"51007710";
		wait for Clk_period;
		Addr <=  "0101110100110";
		Trees_din <= x"b2ffb508";
		wait for Clk_period;
		Addr <=  "0101110100111";
		Trees_din <= x"1afee504";
		wait for Clk_period;
		Addr <=  "0101110101000";
		Trees_din <= x"ffbd2fd5";
		wait for Clk_period;
		Addr <=  "0101110101001";
		Trees_din <= x"004b2fd5";
		wait for Clk_period;
		Addr <=  "0101110101010";
		Trees_din <= x"1efed504";
		wait for Clk_period;
		Addr <=  "0101110101011";
		Trees_din <= x"ffd62fd5";
		wait for Clk_period;
		Addr <=  "0101110101100";
		Trees_din <= x"007b2fd5";
		wait for Clk_period;
		Addr <=  "0101110101101";
		Trees_din <= x"cf000604";
		wait for Clk_period;
		Addr <=  "0101110101110";
		Trees_din <= x"003a2fd5";
		wait for Clk_period;
		Addr <=  "0101110101111";
		Trees_din <= x"ffa32fd5";
		wait for Clk_period;
		Addr <=  "0101110110000";
		Trees_din <= x"91ff4f08";
		wait for Clk_period;
		Addr <=  "0101110110001";
		Trees_din <= x"0bffb604";
		wait for Clk_period;
		Addr <=  "0101110110010";
		Trees_din <= x"00752fd5";
		wait for Clk_period;
		Addr <=  "0101110110011";
		Trees_din <= x"ffeb2fd5";
		wait for Clk_period;
		Addr <=  "0101110110100";
		Trees_din <= x"e2ff4c08";
		wait for Clk_period;
		Addr <=  "0101110110101";
		Trees_din <= x"c5ff0f04";
		wait for Clk_period;
		Addr <=  "0101110110110";
		Trees_din <= x"00042fd5";
		wait for Clk_period;
		Addr <=  "0101110110111";
		Trees_din <= x"ff892fd5";
		wait for Clk_period;
		Addr <=  "0101110111000";
		Trees_din <= x"f3feda04";
		wait for Clk_period;
		Addr <=  "0101110111001";
		Trees_din <= x"00692fd5";
		wait for Clk_period;
		Addr <=  "0101110111010";
		Trees_din <= x"ffe22fd5";
		wait for Clk_period;
		Addr <=  "0101110111011";
		Trees_din <= x"54000f20";
		wait for Clk_period;
		Addr <=  "0101110111100";
		Trees_din <= x"e1ffb310";
		wait for Clk_period;
		Addr <=  "0101110111101";
		Trees_din <= x"32fe3c08";
		wait for Clk_period;
		Addr <=  "0101110111110";
		Trees_din <= x"12ff8e04";
		wait for Clk_period;
		Addr <=  "0101110111111";
		Trees_din <= x"00292fd5";
		wait for Clk_period;
		Addr <=  "0101111000000";
		Trees_din <= x"ff7a2fd5";
		wait for Clk_period;
		Addr <=  "0101111000001";
		Trees_din <= x"33ffce04";
		wait for Clk_period;
		Addr <=  "0101111000010";
		Trees_din <= x"00572fd5";
		wait for Clk_period;
		Addr <=  "0101111000011";
		Trees_din <= x"ffc72fd5";
		wait for Clk_period;
		Addr <=  "0101111000100";
		Trees_din <= x"faffba08";
		wait for Clk_period;
		Addr <=  "0101111000101";
		Trees_din <= x"93ffe504";
		wait for Clk_period;
		Addr <=  "0101111000110";
		Trees_din <= x"fffb2fd5";
		wait for Clk_period;
		Addr <=  "0101111000111";
		Trees_din <= x"ff962fd5";
		wait for Clk_period;
		Addr <=  "0101111001000";
		Trees_din <= x"27004904";
		wait for Clk_period;
		Addr <=  "0101111001001";
		Trees_din <= x"00682fd5";
		wait for Clk_period;
		Addr <=  "0101111001010";
		Trees_din <= x"ffc62fd5";
		wait for Clk_period;
		Addr <=  "0101111001011";
		Trees_din <= x"4cff9510";
		wait for Clk_period;
		Addr <=  "0101111001100";
		Trees_din <= x"1cff4008";
		wait for Clk_period;
		Addr <=  "0101111001101";
		Trees_din <= x"62ff5104";
		wait for Clk_period;
		Addr <=  "0101111001110";
		Trees_din <= x"fffc2fd5";
		wait for Clk_period;
		Addr <=  "0101111001111";
		Trees_din <= x"00322fd5";
		wait for Clk_period;
		Addr <=  "0101111010000";
		Trees_din <= x"ddfec804";
		wait for Clk_period;
		Addr <=  "0101111010001";
		Trees_din <= x"ffbb2fd5";
		wait for Clk_period;
		Addr <=  "0101111010010";
		Trees_din <= x"fff92fd5";
		wait for Clk_period;
		Addr <=  "0101111010011";
		Trees_din <= x"40004b08";
		wait for Clk_period;
		Addr <=  "0101111010100";
		Trees_din <= x"b3ff4104";
		wait for Clk_period;
		Addr <=  "0101111010101";
		Trees_din <= x"ffbe2fd5";
		wait for Clk_period;
		Addr <=  "0101111010110";
		Trees_din <= x"00252fd5";
		wait for Clk_period;
		Addr <=  "0101111010111";
		Trees_din <= x"ff6e2fd5";
		wait for Clk_period;
		Addr <=  "0101111011000";
		Trees_din <= x"6effe510";
		wait for Clk_period;
		Addr <=  "0101111011001";
		Trees_din <= x"9fff3508";
		wait for Clk_period;
		Addr <=  "0101111011010";
		Trees_din <= x"04fff704";
		wait for Clk_period;
		Addr <=  "0101111011011";
		Trees_din <= x"00202fd5";
		wait for Clk_period;
		Addr <=  "0101111011100";
		Trees_din <= x"ff852fd5";
		wait for Clk_period;
		Addr <=  "0101111011101";
		Trees_din <= x"6eff9704";
		wait for Clk_period;
		Addr <=  "0101111011110";
		Trees_din <= x"fffb2fd5";
		wait for Clk_period;
		Addr <=  "0101111011111";
		Trees_din <= x"007b2fd5";
		wait for Clk_period;
		Addr <=  "0101111100000";
		Trees_din <= x"e2ffae20";
		wait for Clk_period;
		Addr <=  "0101111100001";
		Trees_din <= x"56ffed10";
		wait for Clk_period;
		Addr <=  "0101111100010";
		Trees_din <= x"c0ff4d08";
		wait for Clk_period;
		Addr <=  "0101111100011";
		Trees_din <= x"86ff2f04";
		wait for Clk_period;
		Addr <=  "0101111100100";
		Trees_din <= x"ffaf2fd5";
		wait for Clk_period;
		Addr <=  "0101111100101";
		Trees_din <= x"00422fd5";
		wait for Clk_period;
		Addr <=  "0101111100110";
		Trees_din <= x"88ff7504";
		wait for Clk_period;
		Addr <=  "0101111100111";
		Trees_din <= x"00082fd5";
		wait for Clk_period;
		Addr <=  "0101111101000";
		Trees_din <= x"ff772fd5";
		wait for Clk_period;
		Addr <=  "0101111101001";
		Trees_din <= x"cf002008";
		wait for Clk_period;
		Addr <=  "0101111101010";
		Trees_din <= x"1cff9604";
		wait for Clk_period;
		Addr <=  "0101111101011";
		Trees_din <= x"00742fd5";
		wait for Clk_period;
		Addr <=  "0101111101100";
		Trees_din <= x"ffe92fd5";
		wait for Clk_period;
		Addr <=  "0101111101101";
		Trees_din <= x"26004304";
		wait for Clk_period;
		Addr <=  "0101111101110";
		Trees_din <= x"001d2fd5";
		wait for Clk_period;
		Addr <=  "0101111101111";
		Trees_din <= x"ff932fd5";
		wait for Clk_period;
		Addr <=  "0101111110000";
		Trees_din <= x"8e004508";
		wait for Clk_period;
		Addr <=  "0101111110001";
		Trees_din <= x"53ffd004";
		wait for Clk_period;
		Addr <=  "0101111110010";
		Trees_din <= x"00792fd5";
		wait for Clk_period;
		Addr <=  "0101111110011";
		Trees_din <= x"00182fd5";
		wait for Clk_period;
		Addr <=  "0101111110100";
		Trees_din <= x"ffbe2fd5";
		wait for Clk_period;
		Addr <=  "0101111110101";
		Trees_din <= x"d500a264";
		wait for Clk_period;
		Addr <=  "0101111110110";
		Trees_din <= x"67000140";
		wait for Clk_period;
		Addr <=  "0101111110111";
		Trees_din <= x"67ffa420";
		wait for Clk_period;
		Addr <=  "0101111111000";
		Trees_din <= x"31006710";
		wait for Clk_period;
		Addr <=  "0101111111001";
		Trees_din <= x"91ff7508";
		wait for Clk_period;
		Addr <=  "0101111111010";
		Trees_din <= x"c1fe7a04";
		wait for Clk_period;
		Addr <=  "0101111111011";
		Trees_din <= x"002e30b9";
		wait for Clk_period;
		Addr <=  "0101111111100";
		Trees_din <= x"ffe730b9";
		wait for Clk_period;
		Addr <=  "0101111111101";
		Trees_din <= x"81ffa004";
		wait for Clk_period;
		Addr <=  "0101111111110";
		Trees_din <= x"000130b9";
		wait for Clk_period;
		Addr <=  "0101111111111";
		Trees_din <= x"002c30b9";
		wait for Clk_period;
		Addr <=  "0110000000000";
		Trees_din <= x"79ff6308";
		wait for Clk_period;
		Addr <=  "0110000000001";
		Trees_din <= x"f800e404";
		wait for Clk_period;
		Addr <=  "0110000000010";
		Trees_din <= x"ff9b30b9";
		wait for Clk_period;
		Addr <=  "0110000000011";
		Trees_din <= x"003d30b9";
		wait for Clk_period;
		Addr <=  "0110000000100";
		Trees_din <= x"f0ff5c04";
		wait for Clk_period;
		Addr <=  "0110000000101";
		Trees_din <= x"004330b9";
		wait for Clk_period;
		Addr <=  "0110000000110";
		Trees_din <= x"ffdc30b9";
		wait for Clk_period;
		Addr <=  "0110000000111";
		Trees_din <= x"5bffcb10";
		wait for Clk_period;
		Addr <=  "0110000001000";
		Trees_din <= x"62febe08";
		wait for Clk_period;
		Addr <=  "0110000001001";
		Trees_din <= x"55005f04";
		wait for Clk_period;
		Addr <=  "0110000001010";
		Trees_din <= x"007230b9";
		wait for Clk_period;
		Addr <=  "0110000001011";
		Trees_din <= x"ffc030b9";
		wait for Clk_period;
		Addr <=  "0110000001100";
		Trees_din <= x"adff7104";
		wait for Clk_period;
		Addr <=  "0110000001101";
		Trees_din <= x"ffba30b9";
		wait for Clk_period;
		Addr <=  "0110000001110";
		Trees_din <= x"ffef30b9";
		wait for Clk_period;
		Addr <=  "0110000001111";
		Trees_din <= x"a6ff8e08";
		wait for Clk_period;
		Addr <=  "0110000010000";
		Trees_din <= x"c5ff4f04";
		wait for Clk_period;
		Addr <=  "0110000010001";
		Trees_din <= x"008b30b9";
		wait for Clk_period;
		Addr <=  "0110000010010";
		Trees_din <= x"000330b9";
		wait for Clk_period;
		Addr <=  "0110000010011";
		Trees_din <= x"99feca04";
		wait for Clk_period;
		Addr <=  "0110000010100";
		Trees_din <= x"ffa030b9";
		wait for Clk_period;
		Addr <=  "0110000010101";
		Trees_din <= x"002930b9";
		wait for Clk_period;
		Addr <=  "0110000010110";
		Trees_din <= x"89009920";
		wait for Clk_period;
		Addr <=  "0110000010111";
		Trees_din <= x"fbff4c10";
		wait for Clk_period;
		Addr <=  "0110000011000";
		Trees_din <= x"8ffefa08";
		wait for Clk_period;
		Addr <=  "0110000011001";
		Trees_din <= x"a2ff8c04";
		wait for Clk_period;
		Addr <=  "0110000011010";
		Trees_din <= x"ffb530b9";
		wait for Clk_period;
		Addr <=  "0110000011011";
		Trees_din <= x"004830b9";
		wait for Clk_period;
		Addr <=  "0110000011100";
		Trees_din <= x"58ff1d04";
		wait for Clk_period;
		Addr <=  "0110000011101";
		Trees_din <= x"ff7b30b9";
		wait for Clk_period;
		Addr <=  "0110000011110";
		Trees_din <= x"fff930b9";
		wait for Clk_period;
		Addr <=  "0110000011111";
		Trees_din <= x"87ff3c08";
		wait for Clk_period;
		Addr <=  "0110000100000";
		Trees_din <= x"65ff2704";
		wait for Clk_period;
		Addr <=  "0110000100001";
		Trees_din <= x"ff8930b9";
		wait for Clk_period;
		Addr <=  "0110000100010";
		Trees_din <= x"002930b9";
		wait for Clk_period;
		Addr <=  "0110000100011";
		Trees_din <= x"42ff7c04";
		wait for Clk_period;
		Addr <=  "0110000100100";
		Trees_din <= x"008330b9";
		wait for Clk_period;
		Addr <=  "0110000100101";
		Trees_din <= x"002e30b9";
		wait for Clk_period;
		Addr <=  "0110000100110";
		Trees_din <= x"ff9330b9";
		wait for Clk_period;
		Addr <=  "0110000100111";
		Trees_din <= x"78fee008";
		wait for Clk_period;
		Addr <=  "0110000101000";
		Trees_din <= x"03ff7904";
		wait for Clk_period;
		Addr <=  "0110000101001";
		Trees_din <= x"005430b9";
		wait for Clk_period;
		Addr <=  "0110000101010";
		Trees_din <= x"fffd30b9";
		wait for Clk_period;
		Addr <=  "0110000101011";
		Trees_din <= x"24003704";
		wait for Clk_period;
		Addr <=  "0110000101100";
		Trees_din <= x"ff7a30b9";
		wait for Clk_period;
		Addr <=  "0110000101101";
		Trees_din <= x"fff530b9";
		wait for Clk_period;
		Addr <=  "0110000101110";
		Trees_din <= x"a7003c80";
		wait for Clk_period;
		Addr <=  "0110000101111";
		Trees_din <= x"b6ff7240";
		wait for Clk_period;
		Addr <=  "0110000110000";
		Trees_din <= x"24ff9220";
		wait for Clk_period;
		Addr <=  "0110000110001";
		Trees_din <= x"7fff5210";
		wait for Clk_period;
		Addr <=  "0110000110010";
		Trees_din <= x"66ffe908";
		wait for Clk_period;
		Addr <=  "0110000110011";
		Trees_din <= x"afff8b04";
		wait for Clk_period;
		Addr <=  "0110000110100";
		Trees_din <= x"0001324d";
		wait for Clk_period;
		Addr <=  "0110000110101";
		Trees_din <= x"004e324d";
		wait for Clk_period;
		Addr <=  "0110000110110";
		Trees_din <= x"b7ff9704";
		wait for Clk_period;
		Addr <=  "0110000110111";
		Trees_din <= x"ffa8324d";
		wait for Clk_period;
		Addr <=  "0110000111000";
		Trees_din <= x"001e324d";
		wait for Clk_period;
		Addr <=  "0110000111001";
		Trees_din <= x"0d001508";
		wait for Clk_period;
		Addr <=  "0110000111010";
		Trees_din <= x"75ff8e04";
		wait for Clk_period;
		Addr <=  "0110000111011";
		Trees_din <= x"002e324d";
		wait for Clk_period;
		Addr <=  "0110000111100";
		Trees_din <= x"ffc0324d";
		wait for Clk_period;
		Addr <=  "0110000111101";
		Trees_din <= x"e7ff4504";
		wait for Clk_period;
		Addr <=  "0110000111110";
		Trees_din <= x"ffbf324d";
		wait for Clk_period;
		Addr <=  "0110000111111";
		Trees_din <= x"0075324d";
		wait for Clk_period;
		Addr <=  "0110001000000";
		Trees_din <= x"4cfeb310";
		wait for Clk_period;
		Addr <=  "0110001000001";
		Trees_din <= x"5affde08";
		wait for Clk_period;
		Addr <=  "0110001000010";
		Trees_din <= x"3cfef304";
		wait for Clk_period;
		Addr <=  "0110001000011";
		Trees_din <= x"ff9c324d";
		wait for Clk_period;
		Addr <=  "0110001000100";
		Trees_din <= x"ffef324d";
		wait for Clk_period;
		Addr <=  "0110001000101";
		Trees_din <= x"6f002c04";
		wait for Clk_period;
		Addr <=  "0110001000110";
		Trees_din <= x"005d324d";
		wait for Clk_period;
		Addr <=  "0110001000111";
		Trees_din <= x"ffbb324d";
		wait for Clk_period;
		Addr <=  "0110001001000";
		Trees_din <= x"1aff3f08";
		wait for Clk_period;
		Addr <=  "0110001001001";
		Trees_din <= x"e1ff6504";
		wait for Clk_period;
		Addr <=  "0110001001010";
		Trees_din <= x"0038324d";
		wait for Clk_period;
		Addr <=  "0110001001011";
		Trees_din <= x"fff5324d";
		wait for Clk_period;
		Addr <=  "0110001001100";
		Trees_din <= x"adffc304";
		wait for Clk_period;
		Addr <=  "0110001001101";
		Trees_din <= x"004d324d";
		wait for Clk_period;
		Addr <=  "0110001001110";
		Trees_din <= x"fff0324d";
		wait for Clk_period;
		Addr <=  "0110001001111";
		Trees_din <= x"24fffd20";
		wait for Clk_period;
		Addr <=  "0110001010000";
		Trees_din <= x"a0fe3d10";
		wait for Clk_period;
		Addr <=  "0110001010001";
		Trees_din <= x"cbff7d08";
		wait for Clk_period;
		Addr <=  "0110001010010";
		Trees_din <= x"1efff904";
		wait for Clk_period;
		Addr <=  "0110001010011";
		Trees_din <= x"ff7a324d";
		wait for Clk_period;
		Addr <=  "0110001010100";
		Trees_din <= x"0022324d";
		wait for Clk_period;
		Addr <=  "0110001010101";
		Trees_din <= x"a1fe6704";
		wait for Clk_period;
		Addr <=  "0110001010110";
		Trees_din <= x"ffe2324d";
		wait for Clk_period;
		Addr <=  "0110001010111";
		Trees_din <= x"0062324d";
		wait for Clk_period;
		Addr <=  "0110001011000";
		Trees_din <= x"d8ffe908";
		wait for Clk_period;
		Addr <=  "0110001011001";
		Trees_din <= x"e5fec404";
		wait for Clk_period;
		Addr <=  "0110001011010";
		Trees_din <= x"ffe2324d";
		wait for Clk_period;
		Addr <=  "0110001011011";
		Trees_din <= x"0071324d";
		wait for Clk_period;
		Addr <=  "0110001011100";
		Trees_din <= x"ec003b04";
		wait for Clk_period;
		Addr <=  "0110001011101";
		Trees_din <= x"ffcd324d";
		wait for Clk_period;
		Addr <=  "0110001011110";
		Trees_din <= x"0017324d";
		wait for Clk_period;
		Addr <=  "0110001011111";
		Trees_din <= x"a8ff4810";
		wait for Clk_period;
		Addr <=  "0110001100000";
		Trees_din <= x"adff8408";
		wait for Clk_period;
		Addr <=  "0110001100001";
		Trees_din <= x"4dfe7a04";
		wait for Clk_period;
		Addr <=  "0110001100010";
		Trees_din <= x"0060324d";
		wait for Clk_period;
		Addr <=  "0110001100011";
		Trees_din <= x"ffd2324d";
		wait for Clk_period;
		Addr <=  "0110001100100";
		Trees_din <= x"1aff2804";
		wait for Clk_period;
		Addr <=  "0110001100101";
		Trees_din <= x"ff86324d";
		wait for Clk_period;
		Addr <=  "0110001100110";
		Trees_din <= x"0042324d";
		wait for Clk_period;
		Addr <=  "0110001100111";
		Trees_din <= x"2bffaa08";
		wait for Clk_period;
		Addr <=  "0110001101000";
		Trees_din <= x"40001304";
		wait for Clk_period;
		Addr <=  "0110001101001";
		Trees_din <= x"0048324d";
		wait for Clk_period;
		Addr <=  "0110001101010";
		Trees_din <= x"ffd1324d";
		wait for Clk_period;
		Addr <=  "0110001101011";
		Trees_din <= x"de00c504";
		wait for Clk_period;
		Addr <=  "0110001101100";
		Trees_din <= x"007b324d";
		wait for Clk_period;
		Addr <=  "0110001101101";
		Trees_din <= x"ffeb324d";
		wait for Clk_period;
		Addr <=  "0110001101110";
		Trees_din <= x"09fe591c";
		wait for Clk_period;
		Addr <=  "0110001101111";
		Trees_din <= x"95ff1010";
		wait for Clk_period;
		Addr <=  "0110001110000";
		Trees_din <= x"f4ff1c08";
		wait for Clk_period;
		Addr <=  "0110001110001";
		Trees_din <= x"c1febb04";
		wait for Clk_period;
		Addr <=  "0110001110010";
		Trees_din <= x"ff88324d";
		wait for Clk_period;
		Addr <=  "0110001110011";
		Trees_din <= x"0001324d";
		wait for Clk_period;
		Addr <=  "0110001110100";
		Trees_din <= x"b8ff0804";
		wait for Clk_period;
		Addr <=  "0110001110101";
		Trees_din <= x"ffda324d";
		wait for Clk_period;
		Addr <=  "0110001110110";
		Trees_din <= x"005c324d";
		wait for Clk_period;
		Addr <=  "0110001110111";
		Trees_din <= x"d1ff4008";
		wait for Clk_period;
		Addr <=  "0110001111000";
		Trees_din <= x"fcff2b04";
		wait for Clk_period;
		Addr <=  "0110001111001";
		Trees_din <= x"0088324d";
		wait for Clk_period;
		Addr <=  "0110001111010";
		Trees_din <= x"000b324d";
		wait for Clk_period;
		Addr <=  "0110001111011";
		Trees_din <= x"ffca324d";
		wait for Clk_period;
		Addr <=  "0110001111100";
		Trees_din <= x"45ff0818";
		wait for Clk_period;
		Addr <=  "0110001111101";
		Trees_din <= x"b6ff500c";
		wait for Clk_period;
		Addr <=  "0110001111110";
		Trees_din <= x"f202fb08";
		wait for Clk_period;
		Addr <=  "0110001111111";
		Trees_din <= x"8aff7304";
		wait for Clk_period;
		Addr <=  "0110010000000";
		Trees_din <= x"ffcb324d";
		wait for Clk_period;
		Addr <=  "0110010000001";
		Trees_din <= x"ff5a324d";
		wait for Clk_period;
		Addr <=  "0110010000010";
		Trees_din <= x"fff6324d";
		wait for Clk_period;
		Addr <=  "0110010000011";
		Trees_din <= x"32fe6a04";
		wait for Clk_period;
		Addr <=  "0110010000100";
		Trees_din <= x"004c324d";
		wait for Clk_period;
		Addr <=  "0110010000101";
		Trees_din <= x"b3ff4004";
		wait for Clk_period;
		Addr <=  "0110010000110";
		Trees_din <= x"ff97324d";
		wait for Clk_period;
		Addr <=  "0110010000111";
		Trees_din <= x"0022324d";
		wait for Clk_period;
		Addr <=  "0110010001000";
		Trees_din <= x"bdffb908";
		wait for Clk_period;
		Addr <=  "0110010001001";
		Trees_din <= x"c7fedc04";
		wait for Clk_period;
		Addr <=  "0110010001010";
		Trees_din <= x"fff9324d";
		wait for Clk_period;
		Addr <=  "0110010001011";
		Trees_din <= x"006a324d";
		wait for Clk_period;
		Addr <=  "0110010001100";
		Trees_din <= x"d7006008";
		wait for Clk_period;
		Addr <=  "0110010001101";
		Trees_din <= x"44ffc304";
		wait for Clk_period;
		Addr <=  "0110010001110";
		Trees_din <= x"0052324d";
		wait for Clk_period;
		Addr <=  "0110010001111";
		Trees_din <= x"ffca324d";
		wait for Clk_period;
		Addr <=  "0110010010000";
		Trees_din <= x"74ffe204";
		wait for Clk_period;
		Addr <=  "0110010010001";
		Trees_din <= x"ffe1324d";
		wait for Clk_period;
		Addr <=  "0110010010010";
		Trees_din <= x"ff8c324d";
		wait for Clk_period;
		Addr <=  "0110010010011";
		Trees_din <= x"63ffd654";
		wait for Clk_period;
		Addr <=  "0110010010100";
		Trees_din <= x"59008238";
		wait for Clk_period;
		Addr <=  "0110010010101";
		Trees_din <= x"d700f820";
		wait for Clk_period;
		Addr <=  "0110010010110";
		Trees_din <= x"cafdaa10";
		wait for Clk_period;
		Addr <=  "0110010010111";
		Trees_din <= x"17007708";
		wait for Clk_period;
		Addr <=  "0110010011000";
		Trees_din <= x"07ffbc04";
		wait for Clk_period;
		Addr <=  "0110010011001";
		Trees_din <= x"001433c1";
		wait for Clk_period;
		Addr <=  "0110010011010";
		Trees_din <= x"ffac33c1";
		wait for Clk_period;
		Addr <=  "0110010011011";
		Trees_din <= x"3aff7b04";
		wait for Clk_period;
		Addr <=  "0110010011100";
		Trees_din <= x"002033c1";
		wait for Clk_period;
		Addr <=  "0110010011101";
		Trees_din <= x"007e33c1";
		wait for Clk_period;
		Addr <=  "0110010011110";
		Trees_din <= x"76ffb408";
		wait for Clk_period;
		Addr <=  "0110010011111";
		Trees_din <= x"3fffea04";
		wait for Clk_period;
		Addr <=  "0110010100000";
		Trees_din <= x"003433c1";
		wait for Clk_period;
		Addr <=  "0110010100001";
		Trees_din <= x"000733c1";
		wait for Clk_period;
		Addr <=  "0110010100010";
		Trees_din <= x"c9003b04";
		wait for Clk_period;
		Addr <=  "0110010100011";
		Trees_din <= x"000133c1";
		wait for Clk_period;
		Addr <=  "0110010100100";
		Trees_din <= x"ffa833c1";
		wait for Clk_period;
		Addr <=  "0110010100101";
		Trees_din <= x"24ff9e0c";
		wait for Clk_period;
		Addr <=  "0110010100110";
		Trees_din <= x"21ff6504";
		wait for Clk_period;
		Addr <=  "0110010100111";
		Trees_din <= x"ff9933c1";
		wait for Clk_period;
		Addr <=  "0110010101000";
		Trees_din <= x"e3fe6304";
		wait for Clk_period;
		Addr <=  "0110010101001";
		Trees_din <= x"ffa833c1";
		wait for Clk_period;
		Addr <=  "0110010101010";
		Trees_din <= x"005533c1";
		wait for Clk_period;
		Addr <=  "0110010101011";
		Trees_din <= x"cdff4d04";
		wait for Clk_period;
		Addr <=  "0110010101100";
		Trees_din <= x"001133c1";
		wait for Clk_period;
		Addr <=  "0110010101101";
		Trees_din <= x"a8ff7c04";
		wait for Clk_period;
		Addr <=  "0110010101110";
		Trees_din <= x"ff6833c1";
		wait for Clk_period;
		Addr <=  "0110010101111";
		Trees_din <= x"ffce33c1";
		wait for Clk_period;
		Addr <=  "0110010110000";
		Trees_din <= x"26009214";
		wait for Clk_period;
		Addr <=  "0110010110001";
		Trees_din <= x"2cfefe08";
		wait for Clk_period;
		Addr <=  "0110010110010";
		Trees_din <= x"efff9c04";
		wait for Clk_period;
		Addr <=  "0110010110011";
		Trees_din <= x"003b33c1";
		wait for Clk_period;
		Addr <=  "0110010110100";
		Trees_din <= x"ff9d33c1";
		wait for Clk_period;
		Addr <=  "0110010110101";
		Trees_din <= x"6bfeae08";
		wait for Clk_period;
		Addr <=  "0110010110110";
		Trees_din <= x"38ff0304";
		wait for Clk_period;
		Addr <=  "0110010110111";
		Trees_din <= x"ffc333c1";
		wait for Clk_period;
		Addr <=  "0110010111000";
		Trees_din <= x"005833c1";
		wait for Clk_period;
		Addr <=  "0110010111001";
		Trees_din <= x"009033c1";
		wait for Clk_period;
		Addr <=  "0110010111010";
		Trees_din <= x"dcff0004";
		wait for Clk_period;
		Addr <=  "0110010111011";
		Trees_din <= x"002f33c1";
		wait for Clk_period;
		Addr <=  "0110010111100";
		Trees_din <= x"ff8933c1";
		wait for Clk_period;
		Addr <=  "0110010111101";
		Trees_din <= x"6affe13c";
		wait for Clk_period;
		Addr <=  "0110010111110";
		Trees_din <= x"24ffd220";
		wait for Clk_period;
		Addr <=  "0110010111111";
		Trees_din <= x"4afeba10";
		wait for Clk_period;
		Addr <=  "0110011000000";
		Trees_din <= x"a4ffb608";
		wait for Clk_period;
		Addr <=  "0110011000001";
		Trees_din <= x"a4ff7004";
		wait for Clk_period;
		Addr <=  "0110011000010";
		Trees_din <= x"001733c1";
		wait for Clk_period;
		Addr <=  "0110011000011";
		Trees_din <= x"008233c1";
		wait for Clk_period;
		Addr <=  "0110011000100";
		Trees_din <= x"7affd504";
		wait for Clk_period;
		Addr <=  "0110011000101";
		Trees_din <= x"ffa033c1";
		wait for Clk_period;
		Addr <=  "0110011000110";
		Trees_din <= x"000f33c1";
		wait for Clk_period;
		Addr <=  "0110011000111";
		Trees_din <= x"c2ff4008";
		wait for Clk_period;
		Addr <=  "0110011001000";
		Trees_din <= x"d0002c04";
		wait for Clk_period;
		Addr <=  "0110011001001";
		Trees_din <= x"ffbd33c1";
		wait for Clk_period;
		Addr <=  "0110011001010";
		Trees_din <= x"003c33c1";
		wait for Clk_period;
		Addr <=  "0110011001011";
		Trees_din <= x"96ff9504";
		wait for Clk_period;
		Addr <=  "0110011001100";
		Trees_din <= x"ff9833c1";
		wait for Clk_period;
		Addr <=  "0110011001101";
		Trees_din <= x"002633c1";
		wait for Clk_period;
		Addr <=  "0110011001110";
		Trees_din <= x"0bffba0c";
		wait for Clk_period;
		Addr <=  "0110011001111";
		Trees_din <= x"3afecd04";
		wait for Clk_period;
		Addr <=  "0110011010000";
		Trees_din <= x"fffb33c1";
		wait for Clk_period;
		Addr <=  "0110011010001";
		Trees_din <= x"7fffda04";
		wait for Clk_period;
		Addr <=  "0110011010010";
		Trees_din <= x"008e33c1";
		wait for Clk_period;
		Addr <=  "0110011010011";
		Trees_din <= x"001233c1";
		wait for Clk_period;
		Addr <=  "0110011010100";
		Trees_din <= x"82ff5708";
		wait for Clk_period;
		Addr <=  "0110011010101";
		Trees_din <= x"ac001004";
		wait for Clk_period;
		Addr <=  "0110011010110";
		Trees_din <= x"000a33c1";
		wait for Clk_period;
		Addr <=  "0110011010111";
		Trees_din <= x"ff8a33c1";
		wait for Clk_period;
		Addr <=  "0110011011000";
		Trees_din <= x"eaff9104";
		wait for Clk_period;
		Addr <=  "0110011011001";
		Trees_din <= x"ffcf33c1";
		wait for Clk_period;
		Addr <=  "0110011011010";
		Trees_din <= x"006e33c1";
		wait for Clk_period;
		Addr <=  "0110011011011";
		Trees_din <= x"17002318";
		wait for Clk_period;
		Addr <=  "0110011011100";
		Trees_din <= x"3bfee508";
		wait for Clk_period;
		Addr <=  "0110011011101";
		Trees_din <= x"0efe8e04";
		wait for Clk_period;
		Addr <=  "0110011011110";
		Trees_din <= x"ffec33c1";
		wait for Clk_period;
		Addr <=  "0110011011111";
		Trees_din <= x"004433c1";
		wait for Clk_period;
		Addr <=  "0110011100000";
		Trees_din <= x"24000c08";
		wait for Clk_period;
		Addr <=  "0110011100001";
		Trees_din <= x"62fee704";
		wait for Clk_period;
		Addr <=  "0110011100010";
		Trees_din <= x"fff133c1";
		wait for Clk_period;
		Addr <=  "0110011100011";
		Trees_din <= x"ff6f33c1";
		wait for Clk_period;
		Addr <=  "0110011100100";
		Trees_din <= x"e1ffbc04";
		wait for Clk_period;
		Addr <=  "0110011100101";
		Trees_din <= x"ff9c33c1";
		wait for Clk_period;
		Addr <=  "0110011100110";
		Trees_din <= x"003c33c1";
		wait for Clk_period;
		Addr <=  "0110011100111";
		Trees_din <= x"f4ff0e08";
		wait for Clk_period;
		Addr <=  "0110011101000";
		Trees_din <= x"29ffb604";
		wait for Clk_period;
		Addr <=  "0110011101001";
		Trees_din <= x"ff8133c1";
		wait for Clk_period;
		Addr <=  "0110011101010";
		Trees_din <= x"001833c1";
		wait for Clk_period;
		Addr <=  "0110011101011";
		Trees_din <= x"11ff4404";
		wait for Clk_period;
		Addr <=  "0110011101100";
		Trees_din <= x"008833c1";
		wait for Clk_period;
		Addr <=  "0110011101101";
		Trees_din <= x"5cffe904";
		wait for Clk_period;
		Addr <=  "0110011101110";
		Trees_din <= x"003633c1";
		wait for Clk_period;
		Addr <=  "0110011101111";
		Trees_din <= x"ffa733c1";
		wait for Clk_period;
		Addr <=  "0110011110000";
		Trees_din <= x"3100b674";
		wait for Clk_period;
		Addr <=  "0110011110001";
		Trees_din <= x"a6ffaa40";
		wait for Clk_period;
		Addr <=  "0110011110010";
		Trees_din <= x"4fff6120";
		wait for Clk_period;
		Addr <=  "0110011110011";
		Trees_din <= x"a6ff8710";
		wait for Clk_period;
		Addr <=  "0110011110100";
		Trees_din <= x"a6fedc08";
		wait for Clk_period;
		Addr <=  "0110011110101";
		Trees_din <= x"93ff4604";
		wait for Clk_period;
		Addr <=  "0110011110110";
		Trees_din <= x"003334dd";
		wait for Clk_period;
		Addr <=  "0110011110111";
		Trees_din <= x"ffb534dd";
		wait for Clk_period;
		Addr <=  "0110011111000";
		Trees_din <= x"1b001504";
		wait for Clk_period;
		Addr <=  "0110011111001";
		Trees_din <= x"002234dd";
		wait for Clk_period;
		Addr <=  "0110011111010";
		Trees_din <= x"ffe534dd";
		wait for Clk_period;
		Addr <=  "0110011111011";
		Trees_din <= x"37ffea08";
		wait for Clk_period;
		Addr <=  "0110011111100";
		Trees_din <= x"bcfefd04";
		wait for Clk_period;
		Addr <=  "0110011111101";
		Trees_din <= x"ff8b34dd";
		wait for Clk_period;
		Addr <=  "0110011111110";
		Trees_din <= x"fff534dd";
		wait for Clk_period;
		Addr <=  "0110011111111";
		Trees_din <= x"c9ff8f04";
		wait for Clk_period;
		Addr <=  "0110100000000";
		Trees_din <= x"ffd634dd";
		wait for Clk_period;
		Addr <=  "0110100000001";
		Trees_din <= x"005934dd";
		wait for Clk_period;
		Addr <=  "0110100000010";
		Trees_din <= x"91ffee10";
		wait for Clk_period;
		Addr <=  "0110100000011";
		Trees_din <= x"38feef08";
		wait for Clk_period;
		Addr <=  "0110100000100";
		Trees_din <= x"0fff6104";
		wait for Clk_period;
		Addr <=  "0110100000101";
		Trees_din <= x"ffde34dd";
		wait for Clk_period;
		Addr <=  "0110100000110";
		Trees_din <= x"005134dd";
		wait for Clk_period;
		Addr <=  "0110100000111";
		Trees_din <= x"93ff7e04";
		wait for Clk_period;
		Addr <=  "0110100001000";
		Trees_din <= x"fff534dd";
		wait for Clk_period;
		Addr <=  "0110100001001";
		Trees_din <= x"ffca34dd";
		wait for Clk_period;
		Addr <=  "0110100001010";
		Trees_din <= x"b8ff0808";
		wait for Clk_period;
		Addr <=  "0110100001011";
		Trees_din <= x"0dffa404";
		wait for Clk_period;
		Addr <=  "0110100001100";
		Trees_din <= x"ff9b34dd";
		wait for Clk_period;
		Addr <=  "0110100001101";
		Trees_din <= x"000f34dd";
		wait for Clk_period;
		Addr <=  "0110100001110";
		Trees_din <= x"34ffe804";
		wait for Clk_period;
		Addr <=  "0110100001111";
		Trees_din <= x"ffe934dd";
		wait for Clk_period;
		Addr <=  "0110100010000";
		Trees_din <= x"005c34dd";
		wait for Clk_period;
		Addr <=  "0110100010001";
		Trees_din <= x"7dffe814";
		wait for Clk_period;
		Addr <=  "0110100010010";
		Trees_din <= x"51ff0708";
		wait for Clk_period;
		Addr <=  "0110100010011";
		Trees_din <= x"3ffffd04";
		wait for Clk_period;
		Addr <=  "0110100010100";
		Trees_din <= x"001c34dd";
		wait for Clk_period;
		Addr <=  "0110100010101";
		Trees_din <= x"ff8434dd";
		wait for Clk_period;
		Addr <=  "0110100010110";
		Trees_din <= x"d2ff7808";
		wait for Clk_period;
		Addr <=  "0110100010111";
		Trees_din <= x"6ffec204";
		wait for Clk_period;
		Addr <=  "0110100011000";
		Trees_din <= x"ffc134dd";
		wait for Clk_period;
		Addr <=  "0110100011001";
		Trees_din <= x"003e34dd";
		wait for Clk_period;
		Addr <=  "0110100011010";
		Trees_din <= x"ff9d34dd";
		wait for Clk_period;
		Addr <=  "0110100011011";
		Trees_din <= x"6e000c10";
		wait for Clk_period;
		Addr <=  "0110100011100";
		Trees_din <= x"fcfeff08";
		wait for Clk_period;
		Addr <=  "0110100011101";
		Trees_din <= x"15ff7f04";
		wait for Clk_period;
		Addr <=  "0110100011110";
		Trees_din <= x"ff8834dd";
		wait for Clk_period;
		Addr <=  "0110100011111";
		Trees_din <= x"003e34dd";
		wait for Clk_period;
		Addr <=  "0110100100000";
		Trees_din <= x"bd001804";
		wait for Clk_period;
		Addr <=  "0110100100001";
		Trees_din <= x"006a34dd";
		wait for Clk_period;
		Addr <=  "0110100100010";
		Trees_din <= x"ffe034dd";
		wait for Clk_period;
		Addr <=  "0110100100011";
		Trees_din <= x"e7fff608";
		wait for Clk_period;
		Addr <=  "0110100100100";
		Trees_din <= x"86ff5304";
		wait for Clk_period;
		Addr <=  "0110100100101";
		Trees_din <= x"ff9e34dd";
		wait for Clk_period;
		Addr <=  "0110100100110";
		Trees_din <= x"000d34dd";
		wait for Clk_period;
		Addr <=  "0110100100111";
		Trees_din <= x"1fff7f04";
		wait for Clk_period;
		Addr <=  "0110100101000";
		Trees_din <= x"005534dd";
		wait for Clk_period;
		Addr <=  "0110100101001";
		Trees_din <= x"001134dd";
		wait for Clk_period;
		Addr <=  "0110100101010";
		Trees_din <= x"4bfe3004";
		wait for Clk_period;
		Addr <=  "0110100101011";
		Trees_din <= x"003e34dd";
		wait for Clk_period;
		Addr <=  "0110100101100";
		Trees_din <= x"7eff2a14";
		wait for Clk_period;
		Addr <=  "0110100101101";
		Trees_din <= x"54002208";
		wait for Clk_period;
		Addr <=  "0110100101110";
		Trees_din <= x"4cfeed04";
		wait for Clk_period;
		Addr <=  "0110100101111";
		Trees_din <= x"004734dd";
		wait for Clk_period;
		Addr <=  "0110100110000";
		Trees_din <= x"ffa834dd";
		wait for Clk_period;
		Addr <=  "0110100110001";
		Trees_din <= x"be008f08";
		wait for Clk_period;
		Addr <=  "0110100110010";
		Trees_din <= x"cffff804";
		wait for Clk_period;
		Addr <=  "0110100110011";
		Trees_din <= x"ffd234dd";
		wait for Clk_period;
		Addr <=  "0110100110100";
		Trees_din <= x"ff7034dd";
		wait for Clk_period;
		Addr <=  "0110100110101";
		Trees_din <= x"fff234dd";
		wait for Clk_period;
		Addr <=  "0110100110110";
		Trees_din <= x"002a34dd";
		wait for Clk_period;
		Addr <=  "0110100110111";
		Trees_din <= x"d500a26c";
		wait for Clk_period;
		Addr <=  "0110100111000";
		Trees_din <= x"e9fe3f2c";
		wait for Clk_period;
		Addr <=  "0110100111001";
		Trees_din <= x"d3fec814";
		wait for Clk_period;
		Addr <=  "0110100111010";
		Trees_din <= x"32fef60c";
		wait for Clk_period;
		Addr <=  "0110100111011";
		Trees_din <= x"deffa804";
		wait for Clk_period;
		Addr <=  "0110100111100";
		Trees_din <= x"ffcd35c9";
		wait for Clk_period;
		Addr <=  "0110100111101";
		Trees_din <= x"93ff8904";
		wait for Clk_period;
		Addr <=  "0110100111110";
		Trees_din <= x"007f35c9";
		wait for Clk_period;
		Addr <=  "0110100111111";
		Trees_din <= x"ffe835c9";
		wait for Clk_period;
		Addr <=  "0110101000000";
		Trees_din <= x"28ff8704";
		wait for Clk_period;
		Addr <=  "0110101000001";
		Trees_din <= x"ff9b35c9";
		wait for Clk_period;
		Addr <=  "0110101000010";
		Trees_din <= x"002935c9";
		wait for Clk_period;
		Addr <=  "0110101000011";
		Trees_din <= x"7dff4a08";
		wait for Clk_period;
		Addr <=  "0110101000100";
		Trees_din <= x"2cffd504";
		wait for Clk_period;
		Addr <=  "0110101000101";
		Trees_din <= x"006735c9";
		wait for Clk_period;
		Addr <=  "0110101000110";
		Trees_din <= x"ffdf35c9";
		wait for Clk_period;
		Addr <=  "0110101000111";
		Trees_din <= x"9cff8c08";
		wait for Clk_period;
		Addr <=  "0110101001000";
		Trees_din <= x"f4ff3f04";
		wait for Clk_period;
		Addr <=  "0110101001001";
		Trees_din <= x"ff8535c9";
		wait for Clk_period;
		Addr <=  "0110101001010";
		Trees_din <= x"001535c9";
		wait for Clk_period;
		Addr <=  "0110101001011";
		Trees_din <= x"07fffc04";
		wait for Clk_period;
		Addr <=  "0110101001100";
		Trees_din <= x"004035c9";
		wait for Clk_period;
		Addr <=  "0110101001101";
		Trees_din <= x"ffc335c9";
		wait for Clk_period;
		Addr <=  "0110101001110";
		Trees_din <= x"49ffa520";
		wait for Clk_period;
		Addr <=  "0110101001111";
		Trees_din <= x"0bffe310";
		wait for Clk_period;
		Addr <=  "0110101010000";
		Trees_din <= x"f202fe08";
		wait for Clk_period;
		Addr <=  "0110101010001";
		Trees_din <= x"c8ffdb04";
		wait for Clk_period;
		Addr <=  "0110101010010";
		Trees_din <= x"004835c9";
		wait for Clk_period;
		Addr <=  "0110101010011";
		Trees_din <= x"000035c9";
		wait for Clk_period;
		Addr <=  "0110101010100";
		Trees_din <= x"d1ff2504";
		wait for Clk_period;
		Addr <=  "0110101010101";
		Trees_din <= x"ff8235c9";
		wait for Clk_period;
		Addr <=  "0110101010110";
		Trees_din <= x"ffff35c9";
		wait for Clk_period;
		Addr <=  "0110101010111";
		Trees_din <= x"e1ff6d08";
		wait for Clk_period;
		Addr <=  "0110101011000";
		Trees_din <= x"acffd304";
		wait for Clk_period;
		Addr <=  "0110101011001";
		Trees_din <= x"ffad35c9";
		wait for Clk_period;
		Addr <=  "0110101011010";
		Trees_din <= x"005c35c9";
		wait for Clk_period;
		Addr <=  "0110101011011";
		Trees_din <= x"38007104";
		wait for Clk_period;
		Addr <=  "0110101011100";
		Trees_din <= x"ffa935c9";
		wait for Clk_period;
		Addr <=  "0110101011101";
		Trees_din <= x"005635c9";
		wait for Clk_period;
		Addr <=  "0110101011110";
		Trees_din <= x"3dfff810";
		wait for Clk_period;
		Addr <=  "0110101011111";
		Trees_din <= x"20ff6e08";
		wait for Clk_period;
		Addr <=  "0110101100000";
		Trees_din <= x"0efe6804";
		wait for Clk_period;
		Addr <=  "0110101100001";
		Trees_din <= x"ffe835c9";
		wait for Clk_period;
		Addr <=  "0110101100010";
		Trees_din <= x"002c35c9";
		wait for Clk_period;
		Addr <=  "0110101100011";
		Trees_din <= x"45ff4d04";
		wait for Clk_period;
		Addr <=  "0110101100100";
		Trees_din <= x"ffe635c9";
		wait for Clk_period;
		Addr <=  "0110101100101";
		Trees_din <= x"002835c9";
		wait for Clk_period;
		Addr <=  "0110101100110";
		Trees_din <= x"da008308";
		wait for Clk_period;
		Addr <=  "0110101100111";
		Trees_din <= x"96fed004";
		wait for Clk_period;
		Addr <=  "0110101101000";
		Trees_din <= x"ffda35c9";
		wait for Clk_period;
		Addr <=  "0110101101001";
		Trees_din <= x"002735c9";
		wait for Clk_period;
		Addr <=  "0110101101010";
		Trees_din <= x"a7ff0404";
		wait for Clk_period;
		Addr <=  "0110101101011";
		Trees_din <= x"003235c9";
		wait for Clk_period;
		Addr <=  "0110101101100";
		Trees_din <= x"ffa835c9";
		wait for Clk_period;
		Addr <=  "0110101101101";
		Trees_din <= x"78fee004";
		wait for Clk_period;
		Addr <=  "0110101101110";
		Trees_din <= x"002d35c9";
		wait for Clk_period;
		Addr <=  "0110101101111";
		Trees_din <= x"b6ff0004";
		wait for Clk_period;
		Addr <=  "0110101110000";
		Trees_din <= x"ffe435c9";
		wait for Clk_period;
		Addr <=  "0110101110001";
		Trees_din <= x"ff7935c9";
		wait for Clk_period;
		Addr <=  "0110101110010";
		Trees_din <= x"4effff6c";
		wait for Clk_period;
		Addr <=  "0110101110011";
		Trees_din <= x"54002538";
		wait for Clk_period;
		Addr <=  "0110101110100";
		Trees_din <= x"97fe7d18";
		wait for Clk_period;
		Addr <=  "0110101110101";
		Trees_din <= x"0dffbb0c";
		wait for Clk_period;
		Addr <=  "0110101110110";
		Trees_din <= x"57ff3c08";
		wait for Clk_period;
		Addr <=  "0110101110111";
		Trees_din <= x"c2ff2104";
		wait for Clk_period;
		Addr <=  "0110101111000";
		Trees_din <= x"ffee3705";
		wait for Clk_period;
		Addr <=  "0110101111001";
		Trees_din <= x"ff763705";
		wait for Clk_period;
		Addr <=  "0110101111010";
		Trees_din <= x"001b3705";
		wait for Clk_period;
		Addr <=  "0110101111011";
		Trees_din <= x"68feb704";
		wait for Clk_period;
		Addr <=  "0110101111100";
		Trees_din <= x"ffbb3705";
		wait for Clk_period;
		Addr <=  "0110101111101";
		Trees_din <= x"1eff8104";
		wait for Clk_period;
		Addr <=  "0110101111110";
		Trees_din <= x"fff33705";
		wait for Clk_period;
		Addr <=  "0110101111111";
		Trees_din <= x"00743705";
		wait for Clk_period;
		Addr <=  "0110110000000";
		Trees_din <= x"6affc910";
		wait for Clk_period;
		Addr <=  "0110110000001";
		Trees_din <= x"08003108";
		wait for Clk_period;
		Addr <=  "0110110000010";
		Trees_din <= x"3effe604";
		wait for Clk_period;
		Addr <=  "0110110000011";
		Trees_din <= x"00603705";
		wait for Clk_period;
		Addr <=  "0110110000100";
		Trees_din <= x"ffce3705";
		wait for Clk_period;
		Addr <=  "0110110000101";
		Trees_din <= x"e0fed504";
		wait for Clk_period;
		Addr <=  "0110110000110";
		Trees_din <= x"ffe13705";
		wait for Clk_period;
		Addr <=  "0110110000111";
		Trees_din <= x"002d3705";
		wait for Clk_period;
		Addr <=  "0110110001000";
		Trees_din <= x"3eff4a08";
		wait for Clk_period;
		Addr <=  "0110110001001";
		Trees_din <= x"60ff8e04";
		wait for Clk_period;
		Addr <=  "0110110001010";
		Trees_din <= x"00593705";
		wait for Clk_period;
		Addr <=  "0110110001011";
		Trees_din <= x"ffe53705";
		wait for Clk_period;
		Addr <=  "0110110001100";
		Trees_din <= x"45ff0204";
		wait for Clk_period;
		Addr <=  "0110110001101";
		Trees_din <= x"ffba3705";
		wait for Clk_period;
		Addr <=  "0110110001110";
		Trees_din <= x"00123705";
		wait for Clk_period;
		Addr <=  "0110110001111";
		Trees_din <= x"53fff81c";
		wait for Clk_period;
		Addr <=  "0110110010000";
		Trees_din <= x"76002b10";
		wait for Clk_period;
		Addr <=  "0110110010001";
		Trees_din <= x"33ff5a08";
		wait for Clk_period;
		Addr <=  "0110110010010";
		Trees_din <= x"e3fea804";
		wait for Clk_period;
		Addr <=  "0110110010011";
		Trees_din <= x"ffdf3705";
		wait for Clk_period;
		Addr <=  "0110110010100";
		Trees_din <= x"00073705";
		wait for Clk_period;
		Addr <=  "0110110010101";
		Trees_din <= x"8effcb04";
		wait for Clk_period;
		Addr <=  "0110110010110";
		Trees_din <= x"00463705";
		wait for Clk_period;
		Addr <=  "0110110010111";
		Trees_din <= x"000a3705";
		wait for Clk_period;
		Addr <=  "0110110011000";
		Trees_din <= x"57ff8d08";
		wait for Clk_period;
		Addr <=  "0110110011001";
		Trees_din <= x"e8ff6a04";
		wait for Clk_period;
		Addr <=  "0110110011010";
		Trees_din <= x"ff893705";
		wait for Clk_period;
		Addr <=  "0110110011011";
		Trees_din <= x"ffed3705";
		wait for Clk_period;
		Addr <=  "0110110011100";
		Trees_din <= x"00493705";
		wait for Clk_period;
		Addr <=  "0110110011101";
		Trees_din <= x"0dff560c";
		wait for Clk_period;
		Addr <=  "0110110011110";
		Trees_din <= x"c0ff7a08";
		wait for Clk_period;
		Addr <=  "0110110011111";
		Trees_din <= x"e8ff7804";
		wait for Clk_period;
		Addr <=  "0110110100000";
		Trees_din <= x"ffd93705";
		wait for Clk_period;
		Addr <=  "0110110100001";
		Trees_din <= x"00633705";
		wait for Clk_period;
		Addr <=  "0110110100010";
		Trees_din <= x"ffaa3705";
		wait for Clk_period;
		Addr <=  "0110110100011";
		Trees_din <= x"50ffdc08";
		wait for Clk_period;
		Addr <=  "0110110100100";
		Trees_din <= x"56ff1b04";
		wait for Clk_period;
		Addr <=  "0110110100101";
		Trees_din <= x"00073705";
		wait for Clk_period;
		Addr <=  "0110110100110";
		Trees_din <= x"ff843705";
		wait for Clk_period;
		Addr <=  "0110110100111";
		Trees_din <= x"00473705";
		wait for Clk_period;
		Addr <=  "0110110101000";
		Trees_din <= x"bfff7714";
		wait for Clk_period;
		Addr <=  "0110110101001";
		Trees_din <= x"97fe5d04";
		wait for Clk_period;
		Addr <=  "0110110101010";
		Trees_din <= x"00323705";
		wait for Clk_period;
		Addr <=  "0110110101011";
		Trees_din <= x"e4ff540c";
		wait for Clk_period;
		Addr <=  "0110110101100";
		Trees_din <= x"c3ff6304";
		wait for Clk_period;
		Addr <=  "0110110101101";
		Trees_din <= x"fff93705";
		wait for Clk_period;
		Addr <=  "0110110101110";
		Trees_din <= x"14fe8704";
		wait for Clk_period;
		Addr <=  "0110110101111";
		Trees_din <= x"ffe03705";
		wait for Clk_period;
		Addr <=  "0110110110000";
		Trees_din <= x"ff6a3705";
		wait for Clk_period;
		Addr <=  "0110110110001";
		Trees_din <= x"003d3705";
		wait for Clk_period;
		Addr <=  "0110110110010";
		Trees_din <= x"1dfed408";
		wait for Clk_period;
		Addr <=  "0110110110011";
		Trees_din <= x"4afefe04";
		wait for Clk_period;
		Addr <=  "0110110110100";
		Trees_din <= x"fffd3705";
		wait for Clk_period;
		Addr <=  "0110110110101";
		Trees_din <= x"006f3705";
		wait for Clk_period;
		Addr <=  "0110110110110";
		Trees_din <= x"05002610";
		wait for Clk_period;
		Addr <=  "0110110110111";
		Trees_din <= x"51000708";
		wait for Clk_period;
		Addr <=  "0110110111000";
		Trees_din <= x"c6ff4f04";
		wait for Clk_period;
		Addr <=  "0110110111001";
		Trees_din <= x"ffe33705";
		wait for Clk_period;
		Addr <=  "0110110111010";
		Trees_din <= x"00673705";
		wait for Clk_period;
		Addr <=  "0110110111011";
		Trees_din <= x"96ff3a04";
		wait for Clk_period;
		Addr <=  "0110110111100";
		Trees_din <= x"ffa33705";
		wait for Clk_period;
		Addr <=  "0110110111101";
		Trees_din <= x"fff33705";
		wait for Clk_period;
		Addr <=  "0110110111110";
		Trees_din <= x"1effec04";
		wait for Clk_period;
		Addr <=  "0110110111111";
		Trees_din <= x"ff8f3705";
		wait for Clk_period;
		Addr <=  "0110111000000";
		Trees_din <= x"ffeb3705";
		wait for Clk_period;
		Addr <=  "0110111000001";
		Trees_din <= x"59007d70";
		wait for Clk_period;
		Addr <=  "0110111000010";
		Trees_din <= x"05ffea30";
		wait for Clk_period;
		Addr <=  "0110111000011";
		Trees_din <= x"41ff241c";
		wait for Clk_period;
		Addr <=  "0110111000100";
		Trees_din <= x"a9ffdc10";
		wait for Clk_period;
		Addr <=  "0110111000101";
		Trees_din <= x"7d000c08";
		wait for Clk_period;
		Addr <=  "0110111000110";
		Trees_din <= x"2fffbe04";
		wait for Clk_period;
		Addr <=  "0110111000111";
		Trees_din <= x"00793841";
		wait for Clk_period;
		Addr <=  "0110111001000";
		Trees_din <= x"00083841";
		wait for Clk_period;
		Addr <=  "0110111001001";
		Trees_din <= x"35fe9604";
		wait for Clk_period;
		Addr <=  "0110111001010";
		Trees_din <= x"00543841";
		wait for Clk_period;
		Addr <=  "0110111001011";
		Trees_din <= x"ffc33841";
		wait for Clk_period;
		Addr <=  "0110111001100";
		Trees_din <= x"86fed904";
		wait for Clk_period;
		Addr <=  "0110111001101";
		Trees_din <= x"005a3841";
		wait for Clk_period;
		Addr <=  "0110111001110";
		Trees_din <= x"3dffed04";
		wait for Clk_period;
		Addr <=  "0110111001111";
		Trees_din <= x"ff9e3841";
		wait for Clk_period;
		Addr <=  "0110111010000";
		Trees_din <= x"001f3841";
		wait for Clk_period;
		Addr <=  "0110111010001";
		Trees_din <= x"ccff4d08";
		wait for Clk_period;
		Addr <=  "0110111010010";
		Trees_din <= x"ebff4b04";
		wait for Clk_period;
		Addr <=  "0110111010011";
		Trees_din <= x"006e3841";
		wait for Clk_period;
		Addr <=  "0110111010100";
		Trees_din <= x"ffcd3841";
		wait for Clk_period;
		Addr <=  "0110111010101";
		Trees_din <= x"1fff0504";
		wait for Clk_period;
		Addr <=  "0110111010110";
		Trees_din <= x"003f3841";
		wait for Clk_period;
		Addr <=  "0110111010111";
		Trees_din <= x"7c002a04";
		wait for Clk_period;
		Addr <=  "0110111011000";
		Trees_din <= x"ffb53841";
		wait for Clk_period;
		Addr <=  "0110111011001";
		Trees_din <= x"00473841";
		wait for Clk_period;
		Addr <=  "0110111011010";
		Trees_din <= x"3eff9620";
		wait for Clk_period;
		Addr <=  "0110111011011";
		Trees_din <= x"5bffba10";
		wait for Clk_period;
		Addr <=  "0110111011100";
		Trees_din <= x"d9ffe608";
		wait for Clk_period;
		Addr <=  "0110111011101";
		Trees_din <= x"66ffe004";
		wait for Clk_period;
		Addr <=  "0110111011110";
		Trees_din <= x"00133841";
		wait for Clk_period;
		Addr <=  "0110111011111";
		Trees_din <= x"ffe93841";
		wait for Clk_period;
		Addr <=  "0110111100000";
		Trees_din <= x"b3ff4104";
		wait for Clk_period;
		Addr <=  "0110111100001";
		Trees_din <= x"ffc73841";
		wait for Clk_period;
		Addr <=  "0110111100010";
		Trees_din <= x"00063841";
		wait for Clk_period;
		Addr <=  "0110111100011";
		Trees_din <= x"fafef608";
		wait for Clk_period;
		Addr <=  "0110111100100";
		Trees_din <= x"63ff6204";
		wait for Clk_period;
		Addr <=  "0110111100101";
		Trees_din <= x"00153841";
		wait for Clk_period;
		Addr <=  "0110111100110";
		Trees_din <= x"ff923841";
		wait for Clk_period;
		Addr <=  "0110111100111";
		Trees_din <= x"0700cb04";
		wait for Clk_period;
		Addr <=  "0110111101000";
		Trees_din <= x"00473841";
		wait for Clk_period;
		Addr <=  "0110111101001";
		Trees_din <= x"ffcf3841";
		wait for Clk_period;
		Addr <=  "0110111101010";
		Trees_din <= x"d8004410";
		wait for Clk_period;
		Addr <=  "0110111101011";
		Trees_din <= x"e3fed008";
		wait for Clk_period;
		Addr <=  "0110111101100";
		Trees_din <= x"ecff7904";
		wait for Clk_period;
		Addr <=  "0110111101101";
		Trees_din <= x"005c3841";
		wait for Clk_period;
		Addr <=  "0110111101110";
		Trees_din <= x"ffd83841";
		wait for Clk_period;
		Addr <=  "0110111101111";
		Trees_din <= x"e6ffcd04";
		wait for Clk_period;
		Addr <=  "0110111110000";
		Trees_din <= x"fffe3841";
		wait for Clk_period;
		Addr <=  "0110111110001";
		Trees_din <= x"00723841";
		wait for Clk_period;
		Addr <=  "0110111110010";
		Trees_din <= x"43ffb208";
		wait for Clk_period;
		Addr <=  "0110111110011";
		Trees_din <= x"29ffaa04";
		wait for Clk_period;
		Addr <=  "0110111110100";
		Trees_din <= x"ff9c3841";
		wait for Clk_period;
		Addr <=  "0110111110101";
		Trees_din <= x"ffff3841";
		wait for Clk_period;
		Addr <=  "0110111110110";
		Trees_din <= x"20ffc004";
		wait for Clk_period;
		Addr <=  "0110111110111";
		Trees_din <= x"00503841";
		wait for Clk_period;
		Addr <=  "0110111111000";
		Trees_din <= x"ffc43841";
		wait for Clk_period;
		Addr <=  "0110111111001";
		Trees_din <= x"63ffe024";
		wait for Clk_period;
		Addr <=  "0110111111010";
		Trees_din <= x"26006414";
		wait for Clk_period;
		Addr <=  "0110111111011";
		Trees_din <= x"44002f0c";
		wait for Clk_period;
		Addr <=  "0110111111100";
		Trees_din <= x"64fec004";
		wait for Clk_period;
		Addr <=  "0110111111101";
		Trees_din <= x"000b3841";
		wait for Clk_period;
		Addr <=  "0110111111110";
		Trees_din <= x"89003704";
		wait for Clk_period;
		Addr <=  "0110111111111";
		Trees_din <= x"00933841";
		wait for Clk_period;
		Addr <=  "0111000000000";
		Trees_din <= x"00293841";
		wait for Clk_period;
		Addr <=  "0111000000001";
		Trees_din <= x"1fffb804";
		wait for Clk_period;
		Addr <=  "0111000000010";
		Trees_din <= x"004e3841";
		wait for Clk_period;
		Addr <=  "0111000000011";
		Trees_din <= x"ffbe3841";
		wait for Clk_period;
		Addr <=  "0111000000100";
		Trees_din <= x"bfff6708";
		wait for Clk_period;
		Addr <=  "0111000000101";
		Trees_din <= x"f202e404";
		wait for Clk_period;
		Addr <=  "0111000000110";
		Trees_din <= x"00603841";
		wait for Clk_period;
		Addr <=  "0111000000111";
		Trees_din <= x"fff13841";
		wait for Clk_period;
		Addr <=  "0111000001000";
		Trees_din <= x"5a004104";
		wait for Clk_period;
		Addr <=  "0111000001001";
		Trees_din <= x"ff913841";
		wait for Clk_period;
		Addr <=  "0111000001010";
		Trees_din <= x"fff73841";
		wait for Clk_period;
		Addr <=  "0111000001011";
		Trees_din <= x"0a000408";
		wait for Clk_period;
		Addr <=  "0111000001100";
		Trees_din <= x"20ff7204";
		wait for Clk_period;
		Addr <=  "0111000001101";
		Trees_din <= x"ff8f3841";
		wait for Clk_period;
		Addr <=  "0111000001110";
		Trees_din <= x"ffea3841";
		wait for Clk_period;
		Addr <=  "0111000001111";
		Trees_din <= x"00363841";
		wait for Clk_period;
		Addr <=  "0111000010000";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  1
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"08009c80";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"03ffda40";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"86fef720";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"1b001810";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"1eff7808";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"d6005804";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"00a401cd";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"021d01cd";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"d6008904";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"ffe401cd";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"00c201cd";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"3bff6a08";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"b3ff0204";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"01d501cd";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"fff701cd";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"60ff1604";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"ffa401cd";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"039101cd";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"54002710";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"0fffa308";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"5c00f404";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"ff6d01cd";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"00c201cd";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"e4ff5904";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"ffcf01cd";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"015e01cd";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"33fef708";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"47004104";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"005601cd";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"028f01cd";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"7bfed604";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"00a101cd";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"ffc501cd";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"6e006820";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"86fecf10";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"5a008108";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"3afff704";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"029001cd";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"ff8401cd";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"f1ff5204";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"01fb01cd";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"ffdb01cd";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"7bff5d08";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"d3ff5804";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"005a01cd";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"01db01cd";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"18001004";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"ffa301cd";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"011701cd";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"1e001510";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"ceffc008";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"5dff9b04";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"01e901cd";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"008a01cd";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"e1ff9404";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"012d01cd";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"031201cd";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"52feef08";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"13007204";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"ffa401cd";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"030501cd";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"52ffac04";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"ffb501cd";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"016b01cd";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"5cffd73c";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"0700ef20";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"7affda10";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"c7fedf08";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"8b004c04";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"ff5901cd";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"00c201cd";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"be000204";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"ffc001cd";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"016701cd";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"6bfe8508";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"f8006804";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"033301cd";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"fff301cd";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"62ff0204";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"01a101cd";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"ffe401cd";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"8cffcf0c";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"a4ff8b04";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"ff7301cd";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"45ff0204";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"022001cd";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"ff8c01cd";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"0a005908";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"4bfe5804";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"00ca01cd";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"03de01cd";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"01febe04";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"ff9001cd";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"015c01cd";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"77ffee20";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"04ffdd10";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"73fff808";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"60ffcc04";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"ff7101cd";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"00f601cd";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"53ff9d04";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"000001cd";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"02e701cd";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"28fecb08";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"84007f04";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"036801cd";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"008f01cd";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"03ffc204";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"015301cd";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"027801cd";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"dcff0f04";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"01b001cd";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"a4ffe304";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"ff5b01cd";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"008901cd";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"05003278";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"33fefb3c";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"bdffd420";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"62ff4710";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"c1ff0608";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"7bfe7204";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"fffc03a9";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"020403a9";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"43ff4304";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"003c03a9";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"ff7503a9";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"c3ff8308";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"b9feec04";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"ffa403a9";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"025503a9";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"56fef404";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"013b03a9";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"ffcd03a9";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"31004a10";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"5c004d08";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"96feb604";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"00ee03a9";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"ff8a03a9";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"dbfff404";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"ffb503a9";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"016a03a9";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"11ff7808";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"0dff9404";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"023c03a9";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"003003a9";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"ff9303a9";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"7bfef31c";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"86ff6510";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"45ff1c08";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"e9fec304";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"019f03a9";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"007e03a9";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"35fe2304";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"011103a9";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"ff7503a9";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"3100b608";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"0affa704";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"008003a9";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"ff5903a9";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"016f03a9";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"09001e10";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"08007408";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"86fe9204";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"001903a9";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"ff7b03a9";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"62fec504";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"022403a9";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"000203a9";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"6affce08";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"2eff8904";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"009c03a9";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"ff9003a9";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"0cfe9a04";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"001d03a9";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"024903a9";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"3bff2e38";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"e9ff5720";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"11fff310";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"0800dd08";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"53ff7904";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"000d03a9";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"00d103a9";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"21002904";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"019603a9";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"ffd803a9";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"36ffbf08";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"5cff8404";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"008603a9";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"ff5b03a9";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"0b005b04";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"016203a9";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"002e03a9";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"e2ffda10";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"4dfe1e08";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"9fff2604";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"01a303a9";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"ffb503a9";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"a2004204";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"ff6603a9";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"00d303a9";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"08005604";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"ffa703a9";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"01a103a9";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"12ffbf20";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"60ffbe10";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"95fec308";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"1fff6f04";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"ffad03a9";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"017d03a9";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"63ffff04";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"002703a9";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"016403a9";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"d6004508";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"cbff9704";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"017603a9";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"000103a9";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"3fffcf04";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"ffb803a9";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"022103a9";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"54ffc810";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"0f000b08";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"09ffdd04";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"ff6f03a9";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"00ad03a9";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"35fee704";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"001a03a9";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"021d03a9";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"64ff7908";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"83ffb404";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"00f803a9";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"020403a9";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"9ffffe04";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"01f403a9";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"ff8903a9";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"03ff9878";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"aeff2240";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"7aff9c20";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"f2026610";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"20ff7508";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"96001204";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"ff700595";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"007b0595";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"eaff3204";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"01000595";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"ffe30595";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"66ff8108";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"96ff6304";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"01900595";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"ffa40595";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"ebfe6204";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"013a0595";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"ffff0595";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"8e003310";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"26006208";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"09ff9e04";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"ffd00595";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"01070595";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"36ff2b04";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"fff40595";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"00f80595";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"57ff2a08";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"a1ff4d04";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"01de0595";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"00880595";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"0400a604";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"ff8c0595";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"012b0595";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"3bff9c1c";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"99fe450c";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"0afff708";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"03ff3004";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"01e60595";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"00180595";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"ff6e0595";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"6f003e08";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"44005604";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"ff7a0595";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"00030595";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"0dff8804";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"01640595";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"ff890595";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"3effa30c";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"58feed08";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"4aff1104";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"ffe80595";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"01230595";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"ff5b0595";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"2affbf08";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"05000704";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"ff840595";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"00400595";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"67ffdc04";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"02180595";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"00060595";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"28ff1940";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"40003d20";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"8dfeac10";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"3fffac08";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"73000804";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"ff590595";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"009f0595";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"97fe3e04";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"ff7b0595";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"01000595";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"a0feb408";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"ecffbb04";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"ffad0595";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"011f0595";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"faff0904";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"01060595";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"ffc70595";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"a0ff6110";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"36fea808";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"1dff7104";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"ff830595";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"00950595";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"0d007304";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"01780595";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"ff890595";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"0800dd08";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"e7ff7704";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"ff7a0595";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"00c80595";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"6d00eb04";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"01790595";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"00220595";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"54001020";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"aefeee10";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"a2ffdc08";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"3d003704";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"014c0595";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"ffc10595";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"36ff9604";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"ff640595";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"00c90595";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"48fef108";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"00ff8204";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"01b60595";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"ff8b0595";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"52fe9204";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"00680595";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"ff730595";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"d5006a10";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"42ff0708";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"90ffb804";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"01520595";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"ff9a0595";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"12ffe504";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"002a0595";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"009f0595";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"40000a08";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"4eff9d04";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"ff660595";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"00f60595";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"3cff4004";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"02060595";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"006e0595";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"a0ff6570";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"33fef230";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"bd005718";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"9fffd310";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"b3ff8508";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"05002204";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"00430749";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"00e00749";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"baff0c04";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"ff8b0749";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"01660749";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"65ff6804";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"ff530749";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"00ce0749";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"b5fefc10";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"f4ff0b08";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"7dff5904";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"ffd90749";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"011b0749";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"e8febe04";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"00f20749";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"ff740749";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"acffc104";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"003b0749";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"ff580749";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"0700b120";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"1b001310";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"d500a208";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"7bff7f04";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"001f0749";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"ffbf0749";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"e5fe6604";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"ff7c0749";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"015d0749";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"aeff1108";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"39ff9504";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"fff60749";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"01100749";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"eaffa804";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"00560749";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"ff850749";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"74002d10";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"00000508";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"78ff6504";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"01100749";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"00970749";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"68feab04";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"00850749";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"ff5d0749";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"72007508";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"f7002704";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"ffb60749";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"006b0749";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"55006404";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"01820749";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"fff10749";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"54003734";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"0800f020";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"2c001610";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"0f001a08";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"90feee04";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"fff80749";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"ff580749";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"6affdb04";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"ffa30749";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"00d00749";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"5a00ac08";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"49ffff04";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"ff610749";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"006b0749";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"2c004704";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"01d50749";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"ff9c0749";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"fcff5808";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"cbffee04";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"ff690749";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"002a0749";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"83ff2e08";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"e6ff4b04";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"ff930749";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"00210749";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"012d0749";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"3dfffb1c";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"6ffff710";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"5c001808";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"61000604";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"ff9d0749";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"00bb0749";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"f4ff2f04";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"00e20749";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"ff9d0749";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"40ffea04";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"001a0749";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"90ffe504";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"01be0749";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"00330749";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"40007310";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"63ff0808";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"0efe7804";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"011a0749";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"00180749";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"cdff2504";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"00910749";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"ff620749";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"49ffa504";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"ff830749";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"8cffd004";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"00010749";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"01620749";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"54001368";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"f1ffc23c";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"64ff6520";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"08008e10";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"09002e08";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"eafee704";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"00de0915";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"ff9b0915";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"7fff8404";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"ffdc0915";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"00e90915";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"5fff4208";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"b2001504";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"00d90915";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"ffad0915";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"d7010904";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"ff600915";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"007a0915";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"bcff320c";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"2e003408";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"7eff0e04";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"01460915";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"ffb10915";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"ff7e0915";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"11ff3e08";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"2a00be04";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"ff600915";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"002b0915";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"dc001104";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"00c60915";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"ff6f0915";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"8dfe4618";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"93ff3308";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"e0fdcb04";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"001d0915";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"ff620915";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"1300b808";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"c6fe9d04";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"00b80915";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"ff690915";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"7bfef804";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"011e0915";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"00050915";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"44008a0c";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"7c005d08";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"b3ff8a04";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"ff700915";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"00360915";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"00a40915";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"8effdb04";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"ff880915";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"011a0915";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"33fee240";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"3d000320";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"90ff9f10";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"95ff3d08";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"9fffe304";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"010b0915";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"ffae0915";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"33fea804";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"00f20915";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"fff60915";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"1cff4608";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"26007504";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"ff5a0915";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"00830915";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"65febf04";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"ffb90915";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"00c00915";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"28ff0310";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"36ff2908";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"4fff7404";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"ff5b0915";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"008e0915";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"7efee104";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"01000915";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"ffd60915";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"62ff1f08";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"1effdb04";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"00d30915";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"ffa60915";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"f4fe9a04";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"003d0915";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"ff720915";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"05003220";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"da004810";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"64ffc008";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"d3ff7604";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"ffc10915";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"00790915";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"6fff2104";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"010f0915";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"ffc10915";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"05001308";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"20ffc404";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"011a0915";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"ffef0915";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"59001104";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"ff730915";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"007c0915";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"5c001f10";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"8c000e08";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"43ff6f04";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"00400915";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"ffc50915";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"9affa204";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"001d0915";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"00ab0915";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"d6005608";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"ceff8604";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"ffd90915";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"008a0915";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"c8ffc304";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"002f0915";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"00e50915";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"a0ff617c";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"6d005040";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"aeff4520";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"72004810";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"3bff2c08";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"83ffca04";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"ffcf0ac9";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"008d0ac9";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"97fed804";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"fff70ac9";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"006a0ac9";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"90000908";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"04ffca04";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"ffaf0ac9";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"009b0ac9";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"a9ff3904";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"00400ac9";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"ff520ac9";
		wait for Clk_period;
		Addr <=  "0001001010111";
		Trees_din <= x"6e007c10";
		wait for Clk_period;
		Addr <=  "0001001011000";
		Trees_din <= x"f1ff5008";
		wait for Clk_period;
		Addr <=  "0001001011001";
		Trees_din <= x"93ff8c04";
		wait for Clk_period;
		Addr <=  "0001001011010";
		Trees_din <= x"00b90ac9";
		wait for Clk_period;
		Addr <=  "0001001011011";
		Trees_din <= x"ffa30ac9";
		wait for Clk_period;
		Addr <=  "0001001011100";
		Trees_din <= x"fa001b04";
		wait for Clk_period;
		Addr <=  "0001001011101";
		Trees_din <= x"ffa30ac9";
		wait for Clk_period;
		Addr <=  "0001001011110";
		Trees_din <= x"009e0ac9";
		wait for Clk_period;
		Addr <=  "0001001011111";
		Trees_din <= x"03ffdb08";
		wait for Clk_period;
		Addr <=  "0001001100000";
		Trees_din <= x"1800f704";
		wait for Clk_period;
		Addr <=  "0001001100001";
		Trees_din <= x"ffc30ac9";
		wait for Clk_period;
		Addr <=  "0001001100010";
		Trees_din <= x"00c10ac9";
		wait for Clk_period;
		Addr <=  "0001001100011";
		Trees_din <= x"f9fed304";
		wait for Clk_period;
		Addr <=  "0001001100100";
		Trees_din <= x"ffd40ac9";
		wait for Clk_period;
		Addr <=  "0001001100101";
		Trees_din <= x"00e30ac9";
		wait for Clk_period;
		Addr <=  "0001001100110";
		Trees_din <= x"1fffe020";
		wait for Clk_period;
		Addr <=  "0001001100111";
		Trees_din <= x"91ffd210";
		wait for Clk_period;
		Addr <=  "0001001101000";
		Trees_din <= x"8ffe5208";
		wait for Clk_period;
		Addr <=  "0001001101001";
		Trees_din <= x"9ffeeb04";
		wait for Clk_period;
		Addr <=  "0001001101010";
		Trees_din <= x"00e60ac9";
		wait for Clk_period;
		Addr <=  "0001001101011";
		Trees_din <= x"ff930ac9";
		wait for Clk_period;
		Addr <=  "0001001101100";
		Trees_din <= x"f4ff5204";
		wait for Clk_period;
		Addr <=  "0001001101101";
		Trees_din <= x"00a10ac9";
		wait for Clk_period;
		Addr <=  "0001001101110";
		Trees_din <= x"ffc30ac9";
		wait for Clk_period;
		Addr <=  "0001001101111";
		Trees_din <= x"fafff008";
		wait for Clk_period;
		Addr <=  "0001001110000";
		Trees_din <= x"b4fe5b04";
		wait for Clk_period;
		Addr <=  "0001001110001";
		Trees_din <= x"00750ac9";
		wait for Clk_period;
		Addr <=  "0001001110010";
		Trees_din <= x"ff930ac9";
		wait for Clk_period;
		Addr <=  "0001001110011";
		Trees_din <= x"43ff7e04";
		wait for Clk_period;
		Addr <=  "0001001110100";
		Trees_din <= x"01320ac9";
		wait for Clk_period;
		Addr <=  "0001001110101";
		Trees_din <= x"ffaa0ac9";
		wait for Clk_period;
		Addr <=  "0001001110110";
		Trees_din <= x"65001210";
		wait for Clk_period;
		Addr <=  "0001001110111";
		Trees_din <= x"9fff4108";
		wait for Clk_period;
		Addr <=  "0001001111000";
		Trees_din <= x"e3ff5504";
		wait for Clk_period;
		Addr <=  "0001001111001";
		Trees_din <= x"00dc0ac9";
		wait for Clk_period;
		Addr <=  "0001001111010";
		Trees_din <= x"ffcf0ac9";
		wait for Clk_period;
		Addr <=  "0001001111011";
		Trees_din <= x"2bffae04";
		wait for Clk_period;
		Addr <=  "0001001111100";
		Trees_din <= x"00bb0ac9";
		wait for Clk_period;
		Addr <=  "0001001111101";
		Trees_din <= x"00150ac9";
		wait for Clk_period;
		Addr <=  "0001001111110";
		Trees_din <= x"d8005104";
		wait for Clk_period;
		Addr <=  "0001001111111";
		Trees_din <= x"ff5b0ac9";
		wait for Clk_period;
		Addr <=  "0001010000000";
		Trees_din <= x"2aff5a04";
		wait for Clk_period;
		Addr <=  "0001010000001";
		Trees_din <= x"ffec0ac9";
		wait for Clk_period;
		Addr <=  "0001010000010";
		Trees_din <= x"00fd0ac9";
		wait for Clk_period;
		Addr <=  "0001010000011";
		Trees_din <= x"8cffc928";
		wait for Clk_period;
		Addr <=  "0001010000100";
		Trees_din <= x"99fe550c";
		wait for Clk_period;
		Addr <=  "0001010000101";
		Trees_din <= x"5bff6204";
		wait for Clk_period;
		Addr <=  "0001010000110";
		Trees_din <= x"ff850ac9";
		wait for Clk_period;
		Addr <=  "0001010000111";
		Trees_din <= x"96ff2b04";
		wait for Clk_period;
		Addr <=  "0001010001000";
		Trees_din <= x"fff90ac9";
		wait for Clk_period;
		Addr <=  "0001010001001";
		Trees_din <= x"013d0ac9";
		wait for Clk_period;
		Addr <=  "0001010001010";
		Trees_din <= x"e7ffe110";
		wait for Clk_period;
		Addr <=  "0001010001011";
		Trees_din <= x"39003d08";
		wait for Clk_period;
		Addr <=  "0001010001100";
		Trees_din <= x"c1fe0c04";
		wait for Clk_period;
		Addr <=  "0001010001101";
		Trees_din <= x"00410ac9";
		wait for Clk_period;
		Addr <=  "0001010001110";
		Trees_din <= x"ff5f0ac9";
		wait for Clk_period;
		Addr <=  "0001010001111";
		Trees_din <= x"94ff5004";
		wait for Clk_period;
		Addr <=  "0001010010000";
		Trees_din <= x"00b10ac9";
		wait for Clk_period;
		Addr <=  "0001010010001";
		Trees_din <= x"ff8a0ac9";
		wait for Clk_period;
		Addr <=  "0001010010010";
		Trees_din <= x"77fee304";
		wait for Clk_period;
		Addr <=  "0001010010011";
		Trees_din <= x"01160ac9";
		wait for Clk_period;
		Addr <=  "0001010010100";
		Trees_din <= x"75ff8e04";
		wait for Clk_period;
		Addr <=  "0001010010101";
		Trees_din <= x"00740ac9";
		wait for Clk_period;
		Addr <=  "0001010010110";
		Trees_din <= x"ff710ac9";
		wait for Clk_period;
		Addr <=  "0001010010111";
		Trees_din <= x"43ff3e18";
		wait for Clk_period;
		Addr <=  "0001010011000";
		Trees_din <= x"8effc108";
		wait for Clk_period;
		Addr <=  "0001010011001";
		Trees_din <= x"8bff8204";
		wait for Clk_period;
		Addr <=  "0001010011010";
		Trees_din <= x"00760ac9";
		wait for Clk_period;
		Addr <=  "0001010011011";
		Trees_din <= x"ff670ac9";
		wait for Clk_period;
		Addr <=  "0001010011100";
		Trees_din <= x"aeff5308";
		wait for Clk_period;
		Addr <=  "0001010011101";
		Trees_din <= x"7ffebc04";
		wait for Clk_period;
		Addr <=  "0001010011110";
		Trees_din <= x"ffd20ac9";
		wait for Clk_period;
		Addr <=  "0001010011111";
		Trees_din <= x"00fe0ac9";
		wait for Clk_period;
		Addr <=  "0001010100000";
		Trees_din <= x"6fffa804";
		wait for Clk_period;
		Addr <=  "0001010100001";
		Trees_din <= x"ff670ac9";
		wait for Clk_period;
		Addr <=  "0001010100010";
		Trees_din <= x"00a80ac9";
		wait for Clk_period;
		Addr <=  "0001010100011";
		Trees_din <= x"4cff4310";
		wait for Clk_period;
		Addr <=  "0001010100100";
		Trees_din <= x"15ffc508";
		wait for Clk_period;
		Addr <=  "0001010100101";
		Trees_din <= x"2000c104";
		wait for Clk_period;
		Addr <=  "0001010100110";
		Trees_din <= x"ff530ac9";
		wait for Clk_period;
		Addr <=  "0001010100111";
		Trees_din <= x"001a0ac9";
		wait for Clk_period;
		Addr <=  "0001010101000";
		Trees_din <= x"0800bf04";
		wait for Clk_period;
		Addr <=  "0001010101001";
		Trees_din <= x"ffbb0ac9";
		wait for Clk_period;
		Addr <=  "0001010101010";
		Trees_din <= x"00fc0ac9";
		wait for Clk_period;
		Addr <=  "0001010101011";
		Trees_din <= x"0fff6d08";
		wait for Clk_period;
		Addr <=  "0001010101100";
		Trees_din <= x"36ffb704";
		wait for Clk_period;
		Addr <=  "0001010101101";
		Trees_din <= x"ff830ac9";
		wait for Clk_period;
		Addr <=  "0001010101110";
		Trees_din <= x"008e0ac9";
		wait for Clk_period;
		Addr <=  "0001010101111";
		Trees_din <= x"edffbb04";
		wait for Clk_period;
		Addr <=  "0001010110000";
		Trees_din <= x"ffd10ac9";
		wait for Clk_period;
		Addr <=  "0001010110001";
		Trees_din <= x"00d40ac9";
		wait for Clk_period;
		Addr <=  "0001010110010";
		Trees_din <= x"ebff4970";
		wait for Clk_period;
		Addr <=  "0001010110011";
		Trees_din <= x"5fff3c34";
		wait for Clk_period;
		Addr <=  "0001010110100";
		Trees_din <= x"ceffb320";
		wait for Clk_period;
		Addr <=  "0001010110101";
		Trees_din <= x"1effdb10";
		wait for Clk_period;
		Addr <=  "0001010110110";
		Trees_din <= x"05fff908";
		wait for Clk_period;
		Addr <=  "0001010110111";
		Trees_din <= x"7bfef204";
		wait for Clk_period;
		Addr <=  "0001010111000";
		Trees_din <= x"004a0c2d";
		wait for Clk_period;
		Addr <=  "0001010111001";
		Trees_din <= x"ff7d0c2d";
		wait for Clk_period;
		Addr <=  "0001010111010";
		Trees_din <= x"00ff9a04";
		wait for Clk_period;
		Addr <=  "0001010111011";
		Trees_din <= x"00830c2d";
		wait for Clk_period;
		Addr <=  "0001010111100";
		Trees_din <= x"00030c2d";
		wait for Clk_period;
		Addr <=  "0001010111101";
		Trees_din <= x"22007008";
		wait for Clk_period;
		Addr <=  "0001010111110";
		Trees_din <= x"e9fe5904";
		wait for Clk_period;
		Addr <=  "0001010111111";
		Trees_din <= x"00670c2d";
		wait for Clk_period;
		Addr <=  "0001011000000";
		Trees_din <= x"ff900c2d";
		wait for Clk_period;
		Addr <=  "0001011000001";
		Trees_din <= x"0eff5f04";
		wait for Clk_period;
		Addr <=  "0001011000010";
		Trees_din <= x"00070c2d";
		wait for Clk_period;
		Addr <=  "0001011000011";
		Trees_din <= x"012e0c2d";
		wait for Clk_period;
		Addr <=  "0001011000100";
		Trees_din <= x"6dffa004";
		wait for Clk_period;
		Addr <=  "0001011000101";
		Trees_din <= x"ff6a0c2d";
		wait for Clk_period;
		Addr <=  "0001011000110";
		Trees_din <= x"6e000908";
		wait for Clk_period;
		Addr <=  "0001011000111";
		Trees_din <= x"06ff3b04";
		wait for Clk_period;
		Addr <=  "0001011001000";
		Trees_din <= x"00a20c2d";
		wait for Clk_period;
		Addr <=  "0001011001001";
		Trees_din <= x"000c0c2d";
		wait for Clk_period;
		Addr <=  "0001011001010";
		Trees_din <= x"2affbd04";
		wait for Clk_period;
		Addr <=  "0001011001011";
		Trees_din <= x"00620c2d";
		wait for Clk_period;
		Addr <=  "0001011001100";
		Trees_din <= x"00b30c2d";
		wait for Clk_period;
		Addr <=  "0001011001101";
		Trees_din <= x"03ff121c";
		wait for Clk_period;
		Addr <=  "0001011001110";
		Trees_din <= x"6effe610";
		wait for Clk_period;
		Addr <=  "0001011001111";
		Trees_din <= x"06ff4808";
		wait for Clk_period;
		Addr <=  "0001011010000";
		Trees_din <= x"21ffc704";
		wait for Clk_period;
		Addr <=  "0001011010001";
		Trees_din <= x"01620c2d";
		wait for Clk_period;
		Addr <=  "0001011010010";
		Trees_din <= x"ff980c2d";
		wait for Clk_period;
		Addr <=  "0001011010011";
		Trees_din <= x"b6ffbd04";
		wait for Clk_period;
		Addr <=  "0001011010100";
		Trees_din <= x"ff5f0c2d";
		wait for Clk_period;
		Addr <=  "0001011010101";
		Trees_din <= x"00a20c2d";
		wait for Clk_period;
		Addr <=  "0001011010110";
		Trees_din <= x"a6fe8704";
		wait for Clk_period;
		Addr <=  "0001011010111";
		Trees_din <= x"006b0c2d";
		wait for Clk_period;
		Addr <=  "0001011011000";
		Trees_din <= x"8fffa104";
		wait for Clk_period;
		Addr <=  "0001011011001";
		Trees_din <= x"ff510c2d";
		wait for Clk_period;
		Addr <=  "0001011011010";
		Trees_din <= x"002b0c2d";
		wait for Clk_period;
		Addr <=  "0001011011011";
		Trees_din <= x"7aff9c10";
		wait for Clk_period;
		Addr <=  "0001011011100";
		Trees_din <= x"d600ac08";
		wait for Clk_period;
		Addr <=  "0001011011101";
		Trees_din <= x"d2ff9304";
		wait for Clk_period;
		Addr <=  "0001011011110";
		Trees_din <= x"ffde0c2d";
		wait for Clk_period;
		Addr <=  "0001011011111";
		Trees_din <= x"00f40c2d";
		wait for Clk_period;
		Addr <=  "0001011100000";
		Trees_din <= x"36ff1604";
		wait for Clk_period;
		Addr <=  "0001011100001";
		Trees_din <= x"ffc10c2d";
		wait for Clk_period;
		Addr <=  "0001011100010";
		Trees_din <= x"009a0c2d";
		wait for Clk_period;
		Addr <=  "0001011100011";
		Trees_din <= x"0fff1808";
		wait for Clk_period;
		Addr <=  "0001011100100";
		Trees_din <= x"5effe704";
		wait for Clk_period;
		Addr <=  "0001011100101";
		Trees_din <= x"ff7d0c2d";
		wait for Clk_period;
		Addr <=  "0001011100110";
		Trees_din <= x"005e0c2d";
		wait for Clk_period;
		Addr <=  "0001011100111";
		Trees_din <= x"a1ff9804";
		wait for Clk_period;
		Addr <=  "0001011101000";
		Trees_din <= x"00630c2d";
		wait for Clk_period;
		Addr <=  "0001011101001";
		Trees_din <= x"ffa70c2d";
		wait for Clk_period;
		Addr <=  "0001011101010";
		Trees_din <= x"6f005e3c";
		wait for Clk_period;
		Addr <=  "0001011101011";
		Trees_din <= x"62ff5320";
		wait for Clk_period;
		Addr <=  "0001011101100";
		Trees_din <= x"d3fed510";
		wait for Clk_period;
		Addr <=  "0001011101101";
		Trees_din <= x"94008308";
		wait for Clk_period;
		Addr <=  "0001011101110";
		Trees_din <= x"19ff9404";
		wait for Clk_period;
		Addr <=  "0001011101111";
		Trees_din <= x"ff770c2d";
		wait for Clk_period;
		Addr <=  "0001011110000";
		Trees_din <= x"00650c2d";
		wait for Clk_period;
		Addr <=  "0001011110001";
		Trees_din <= x"89ffd604";
		wait for Clk_period;
		Addr <=  "0001011110010";
		Trees_din <= x"00c70c2d";
		wait for Clk_period;
		Addr <=  "0001011110011";
		Trees_din <= x"ffa50c2d";
		wait for Clk_period;
		Addr <=  "0001011110100";
		Trees_din <= x"02fe8b08";
		wait for Clk_period;
		Addr <=  "0001011110101";
		Trees_din <= x"f5ffc704";
		wait for Clk_period;
		Addr <=  "0001011110110";
		Trees_din <= x"00040c2d";
		wait for Clk_period;
		Addr <=  "0001011110111";
		Trees_din <= x"ff630c2d";
		wait for Clk_period;
		Addr <=  "0001011111000";
		Trees_din <= x"ac001304";
		wait for Clk_period;
		Addr <=  "0001011111001";
		Trees_din <= x"00d70c2d";
		wait for Clk_period;
		Addr <=  "0001011111010";
		Trees_din <= x"001b0c2d";
		wait for Clk_period;
		Addr <=  "0001011111011";
		Trees_din <= x"38003a10";
		wait for Clk_period;
		Addr <=  "0001011111100";
		Trees_din <= x"39fec108";
		wait for Clk_period;
		Addr <=  "0001011111101";
		Trees_din <= x"2cffc204";
		wait for Clk_period;
		Addr <=  "0001011111110";
		Trees_din <= x"ff870c2d";
		wait for Clk_period;
		Addr <=  "0001011111111";
		Trees_din <= x"011f0c2d";
		wait for Clk_period;
		Addr <=  "0001100000000";
		Trees_din <= x"6d00b004";
		wait for Clk_period;
		Addr <=  "0001100000001";
		Trees_din <= x"ff660c2d";
		wait for Clk_period;
		Addr <=  "0001100000010";
		Trees_din <= x"00530c2d";
		wait for Clk_period;
		Addr <=  "0001100000011";
		Trees_din <= x"95fef908";
		wait for Clk_period;
		Addr <=  "0001100000100";
		Trees_din <= x"a9ff3304";
		wait for Clk_period;
		Addr <=  "0001100000101";
		Trees_din <= x"00420c2d";
		wait for Clk_period;
		Addr <=  "0001100000110";
		Trees_din <= x"015a0c2d";
		wait for Clk_period;
		Addr <=  "0001100000111";
		Trees_din <= x"ff880c2d";
		wait for Clk_period;
		Addr <=  "0001100001000";
		Trees_din <= x"46ff0004";
		wait for Clk_period;
		Addr <=  "0001100001001";
		Trees_din <= x"003c0c2d";
		wait for Clk_period;
		Addr <=  "0001100001010";
		Trees_din <= x"01470c2d";
		wait for Clk_period;
		Addr <=  "0001100001011";
		Trees_din <= x"43ffa77c";
		wait for Clk_period;
		Addr <=  "0001100001100";
		Trees_din <= x"8cff6440";
		wait for Clk_period;
		Addr <=  "0001100001101";
		Trees_din <= x"36ff5420";
		wait for Clk_period;
		Addr <=  "0001100001110";
		Trees_din <= x"b5fe1810";
		wait for Clk_period;
		Addr <=  "0001100001111";
		Trees_din <= x"9cff3808";
		wait for Clk_period;
		Addr <=  "0001100010000";
		Trees_din <= x"ac002404";
		wait for Clk_period;
		Addr <=  "0001100010001";
		Trees_din <= x"01430de9";
		wait for Clk_period;
		Addr <=  "0001100010010";
		Trees_din <= x"000d0de9";
		wait for Clk_period;
		Addr <=  "0001100010011";
		Trees_din <= x"55ffb204";
		wait for Clk_period;
		Addr <=  "0001100010100";
		Trees_din <= x"00770de9";
		wait for Clk_period;
		Addr <=  "0001100010101";
		Trees_din <= x"ff7d0de9";
		wait for Clk_period;
		Addr <=  "0001100010110";
		Trees_din <= x"be008a08";
		wait for Clk_period;
		Addr <=  "0001100010111";
		Trees_din <= x"b3ff9f04";
		wait for Clk_period;
		Addr <=  "0001100011000";
		Trees_din <= x"ffa50de9";
		wait for Clk_period;
		Addr <=  "0001100011001";
		Trees_din <= x"00a20de9";
		wait for Clk_period;
		Addr <=  "0001100011010";
		Trees_din <= x"80ff7404";
		wait for Clk_period;
		Addr <=  "0001100011011";
		Trees_din <= x"00f00de9";
		wait for Clk_period;
		Addr <=  "0001100011100";
		Trees_din <= x"ffcb0de9";
		wait for Clk_period;
		Addr <=  "0001100011101";
		Trees_din <= x"87ff5f10";
		wait for Clk_period;
		Addr <=  "0001100011110";
		Trees_din <= x"29ff4808";
		wait for Clk_period;
		Addr <=  "0001100011111";
		Trees_din <= x"08ffc304";
		wait for Clk_period;
		Addr <=  "0001100100000";
		Trees_din <= x"ff820de9";
		wait for Clk_period;
		Addr <=  "0001100100001";
		Trees_din <= x"01050de9";
		wait for Clk_period;
		Addr <=  "0001100100010";
		Trees_din <= x"cc003b04";
		wait for Clk_period;
		Addr <=  "0001100100011";
		Trees_din <= x"ffdf0de9";
		wait for Clk_period;
		Addr <=  "0001100100100";
		Trees_din <= x"00c60de9";
		wait for Clk_period;
		Addr <=  "0001100100101";
		Trees_din <= x"5dff9208";
		wait for Clk_period;
		Addr <=  "0001100100110";
		Trees_din <= x"ceff9c04";
		wait for Clk_period;
		Addr <=  "0001100100111";
		Trees_din <= x"ffb50de9";
		wait for Clk_period;
		Addr <=  "0001100101000";
		Trees_din <= x"00d10de9";
		wait for Clk_period;
		Addr <=  "0001100101001";
		Trees_din <= x"b3ff9004";
		wait for Clk_period;
		Addr <=  "0001100101010";
		Trees_din <= x"ffa90de9";
		wait for Clk_period;
		Addr <=  "0001100101011";
		Trees_din <= x"00800de9";
		wait for Clk_period;
		Addr <=  "0001100101100";
		Trees_din <= x"86feff20";
		wait for Clk_period;
		Addr <=  "0001100101101";
		Trees_din <= x"5c002c10";
		wait for Clk_period;
		Addr <=  "0001100101110";
		Trees_din <= x"40003d08";
		wait for Clk_period;
		Addr <=  "0001100101111";
		Trees_din <= x"48fff904";
		wait for Clk_period;
		Addr <=  "0001100110000";
		Trees_din <= x"00480de9";
		wait for Clk_period;
		Addr <=  "0001100110001";
		Trees_din <= x"ffcc0de9";
		wait for Clk_period;
		Addr <=  "0001100110010";
		Trees_din <= x"db007204";
		wait for Clk_period;
		Addr <=  "0001100110011";
		Trees_din <= x"00c20de9";
		wait for Clk_period;
		Addr <=  "0001100110100";
		Trees_din <= x"ffee0de9";
		wait for Clk_period;
		Addr <=  "0001100110101";
		Trees_din <= x"1dfe1d08";
		wait for Clk_period;
		Addr <=  "0001100110110";
		Trees_din <= x"65ff1b04";
		wait for Clk_period;
		Addr <=  "0001100110111";
		Trees_din <= x"00310de9";
		wait for Clk_period;
		Addr <=  "0001100111000";
		Trees_din <= x"ff6e0de9";
		wait for Clk_period;
		Addr <=  "0001100111001";
		Trees_din <= x"74002704";
		wait for Clk_period;
		Addr <=  "0001100111010";
		Trees_din <= x"00ba0de9";
		wait for Clk_period;
		Addr <=  "0001100111011";
		Trees_din <= x"00470de9";
		wait for Clk_period;
		Addr <=  "0001100111100";
		Trees_din <= x"6f003210";
		wait for Clk_period;
		Addr <=  "0001100111101";
		Trees_din <= x"aefecb08";
		wait for Clk_period;
		Addr <=  "0001100111110";
		Trees_din <= x"c3002804";
		wait for Clk_period;
		Addr <=  "0001100111111";
		Trees_din <= x"00340de9";
		wait for Clk_period;
		Addr <=  "0001101000000";
		Trees_din <= x"00ab0de9";
		wait for Clk_period;
		Addr <=  "0001101000001";
		Trees_din <= x"34000804";
		wait for Clk_period;
		Addr <=  "0001101000010";
		Trees_din <= x"ffcc0de9";
		wait for Clk_period;
		Addr <=  "0001101000011";
		Trees_din <= x"002c0de9";
		wait for Clk_period;
		Addr <=  "0001101000100";
		Trees_din <= x"92ffdb08";
		wait for Clk_period;
		Addr <=  "0001101000101";
		Trees_din <= x"e6ff6404";
		wait for Clk_period;
		Addr <=  "0001101000110";
		Trees_din <= x"ffb70de9";
		wait for Clk_period;
		Addr <=  "0001101000111";
		Trees_din <= x"00ed0de9";
		wait for Clk_period;
		Addr <=  "0001101001000";
		Trees_din <= x"ff7e0de9";
		wait for Clk_period;
		Addr <=  "0001101001001";
		Trees_din <= x"31005234";
		wait for Clk_period;
		Addr <=  "0001101001010";
		Trees_din <= x"44008a20";
		wait for Clk_period;
		Addr <=  "0001101001011";
		Trees_din <= x"24ffb810";
		wait for Clk_period;
		Addr <=  "0001101001100";
		Trees_din <= x"ecff9b08";
		wait for Clk_period;
		Addr <=  "0001101001101";
		Trees_din <= x"f1ffc104";
		wait for Clk_period;
		Addr <=  "0001101001110";
		Trees_din <= x"00ba0de9";
		wait for Clk_period;
		Addr <=  "0001101001111";
		Trees_din <= x"ff9b0de9";
		wait for Clk_period;
		Addr <=  "0001101010000";
		Trees_din <= x"c9ffd604";
		wait for Clk_period;
		Addr <=  "0001101010001";
		Trees_din <= x"ff9e0de9";
		wait for Clk_period;
		Addr <=  "0001101010010";
		Trees_din <= x"001e0de9";
		wait for Clk_period;
		Addr <=  "0001101010011";
		Trees_din <= x"1b004c08";
		wait for Clk_period;
		Addr <=  "0001101010100";
		Trees_din <= x"79fed104";
		wait for Clk_period;
		Addr <=  "0001101010101";
		Trees_din <= x"003f0de9";
		wait for Clk_period;
		Addr <=  "0001101010110";
		Trees_din <= x"ff7d0de9";
		wait for Clk_period;
		Addr <=  "0001101010111";
		Trees_din <= x"99ff0204";
		wait for Clk_period;
		Addr <=  "0001101011000";
		Trees_din <= x"00c30de9";
		wait for Clk_period;
		Addr <=  "0001101011001";
		Trees_din <= x"ff7a0de9";
		wait for Clk_period;
		Addr <=  "0001101011010";
		Trees_din <= x"8affe910";
		wait for Clk_period;
		Addr <=  "0001101011011";
		Trees_din <= x"e1ff8308";
		wait for Clk_period;
		Addr <=  "0001101011100";
		Trees_din <= x"7dffd304";
		wait for Clk_period;
		Addr <=  "0001101011101";
		Trees_din <= x"ff9a0de9";
		wait for Clk_period;
		Addr <=  "0001101011110";
		Trees_din <= x"00130de9";
		wait for Clk_period;
		Addr <=  "0001101011111";
		Trees_din <= x"8cff4004";
		wait for Clk_period;
		Addr <=  "0001101100000";
		Trees_din <= x"ffee0de9";
		wait for Clk_period;
		Addr <=  "0001101100001";
		Trees_din <= x"01310de9";
		wait for Clk_period;
		Addr <=  "0001101100010";
		Trees_din <= x"ff6b0de9";
		wait for Clk_period;
		Addr <=  "0001101100011";
		Trees_din <= x"5bffa220";
		wait for Clk_period;
		Addr <=  "0001101100100";
		Trees_din <= x"a0ff7010";
		wait for Clk_period;
		Addr <=  "0001101100101";
		Trees_din <= x"a9ff9008";
		wait for Clk_period;
		Addr <=  "0001101100110";
		Trees_din <= x"5e003104";
		wait for Clk_period;
		Addr <=  "0001101100111";
		Trees_din <= x"010c0de9";
		wait for Clk_period;
		Addr <=  "0001101101000";
		Trees_din <= x"ffe70de9";
		wait for Clk_period;
		Addr <=  "0001101101001";
		Trees_din <= x"7dffaa04";
		wait for Clk_period;
		Addr <=  "0001101101010";
		Trees_din <= x"ff880de9";
		wait for Clk_period;
		Addr <=  "0001101101011";
		Trees_din <= x"009e0de9";
		wait for Clk_period;
		Addr <=  "0001101101100";
		Trees_din <= x"ceffb708";
		wait for Clk_period;
		Addr <=  "0001101101101";
		Trees_din <= x"68fe4104";
		wait for Clk_period;
		Addr <=  "0001101101110";
		Trees_din <= x"fff80de9";
		wait for Clk_period;
		Addr <=  "0001101101111";
		Trees_din <= x"ff710de9";
		wait for Clk_period;
		Addr <=  "0001101110000";
		Trees_din <= x"04009a04";
		wait for Clk_period;
		Addr <=  "0001101110001";
		Trees_din <= x"00080de9";
		wait for Clk_period;
		Addr <=  "0001101110010";
		Trees_din <= x"00810de9";
		wait for Clk_period;
		Addr <=  "0001101110011";
		Trees_din <= x"84ff4608";
		wait for Clk_period;
		Addr <=  "0001101110100";
		Trees_din <= x"11ff3604";
		wait for Clk_period;
		Addr <=  "0001101110101";
		Trees_din <= x"ffe80de9";
		wait for Clk_period;
		Addr <=  "0001101110110";
		Trees_din <= x"00c80de9";
		wait for Clk_period;
		Addr <=  "0001101110111";
		Trees_din <= x"41fe9304";
		wait for Clk_period;
		Addr <=  "0001101111000";
		Trees_din <= x"00120de9";
		wait for Clk_period;
		Addr <=  "0001101111001";
		Trees_din <= x"ff5c0de9";
		wait for Clk_period;
		Addr <=  "0001101111010";
		Trees_din <= x"05003270";
		wait for Clk_period;
		Addr <=  "0001101111011";
		Trees_din <= x"45ff1c3c";
		wait for Clk_period;
		Addr <=  "0001101111100";
		Trees_din <= x"61ff5e1c";
		wait for Clk_period;
		Addr <=  "0001101111101";
		Trees_din <= x"33feaa0c";
		wait for Clk_period;
		Addr <=  "0001101111110";
		Trees_din <= x"80ff3804";
		wait for Clk_period;
		Addr <=  "0001101111111";
		Trees_din <= x"ff760fc5";
		wait for Clk_period;
		Addr <=  "0001110000000";
		Trees_din <= x"54000004";
		wait for Clk_period;
		Addr <=  "0001110000001";
		Trees_din <= x"ff880fc5";
		wait for Clk_period;
		Addr <=  "0001110000010";
		Trees_din <= x"00ad0fc5";
		wait for Clk_period;
		Addr <=  "0001110000011";
		Trees_din <= x"83ff3208";
		wait for Clk_period;
		Addr <=  "0001110000100";
		Trees_din <= x"6afeca04";
		wait for Clk_period;
		Addr <=  "0001110000101";
		Trees_din <= x"009d0fc5";
		wait for Clk_period;
		Addr <=  "0001110000110";
		Trees_din <= x"ff8a0fc5";
		wait for Clk_period;
		Addr <=  "0001110000111";
		Trees_din <= x"1300ac04";
		wait for Clk_period;
		Addr <=  "0001110001000";
		Trees_din <= x"ffa90fc5";
		wait for Clk_period;
		Addr <=  "0001110001001";
		Trees_din <= x"006d0fc5";
		wait for Clk_period;
		Addr <=  "0001110001010";
		Trees_din <= x"20ff2e10";
		wait for Clk_period;
		Addr <=  "0001110001011";
		Trees_din <= x"64ff9e08";
		wait for Clk_period;
		Addr <=  "0001110001100";
		Trees_din <= x"e800a604";
		wait for Clk_period;
		Addr <=  "0001110001101";
		Trees_din <= x"ff7a0fc5";
		wait for Clk_period;
		Addr <=  "0001110001110";
		Trees_din <= x"00b90fc5";
		wait for Clk_period;
		Addr <=  "0001110001111";
		Trees_din <= x"3afeed04";
		wait for Clk_period;
		Addr <=  "0001110010000";
		Trees_din <= x"012c0fc5";
		wait for Clk_period;
		Addr <=  "0001110010001";
		Trees_din <= x"ffd90fc5";
		wait for Clk_period;
		Addr <=  "0001110010010";
		Trees_din <= x"6bfeb908";
		wait for Clk_period;
		Addr <=  "0001110010011";
		Trees_din <= x"96ff7a04";
		wait for Clk_period;
		Addr <=  "0001110010100";
		Trees_din <= x"00d70fc5";
		wait for Clk_period;
		Addr <=  "0001110010101";
		Trees_din <= x"00080fc5";
		wait for Clk_period;
		Addr <=  "0001110010110";
		Trees_din <= x"da004804";
		wait for Clk_period;
		Addr <=  "0001110010111";
		Trees_din <= x"fffc0fc5";
		wait for Clk_period;
		Addr <=  "0001110011000";
		Trees_din <= x"00790fc5";
		wait for Clk_period;
		Addr <=  "0001110011001";
		Trees_din <= x"31ffc714";
		wait for Clk_period;
		Addr <=  "0001110011010";
		Trees_din <= x"79006910";
		wait for Clk_period;
		Addr <=  "0001110011011";
		Trees_din <= x"b3ff8e08";
		wait for Clk_period;
		Addr <=  "0001110011100";
		Trees_din <= x"96fe7a04";
		wait for Clk_period;
		Addr <=  "0001110011101";
		Trees_din <= x"00710fc5";
		wait for Clk_period;
		Addr <=  "0001110011110";
		Trees_din <= x"ff700fc5";
		wait for Clk_period;
		Addr <=  "0001110011111";
		Trees_din <= x"33feef04";
		wait for Clk_period;
		Addr <=  "0001110100000";
		Trees_din <= x"00c30fc5";
		wait for Clk_period;
		Addr <=  "0001110100001";
		Trees_din <= x"ffa10fc5";
		wait for Clk_period;
		Addr <=  "0001110100010";
		Trees_din <= x"01340fc5";
		wait for Clk_period;
		Addr <=  "0001110100011";
		Trees_din <= x"bcfebf10";
		wait for Clk_period;
		Addr <=  "0001110100100";
		Trees_din <= x"10000208";
		wait for Clk_period;
		Addr <=  "0001110100101";
		Trees_din <= x"82ffca04";
		wait for Clk_period;
		Addr <=  "0001110100110";
		Trees_din <= x"01020fc5";
		wait for Clk_period;
		Addr <=  "0001110100111";
		Trees_din <= x"ffde0fc5";
		wait for Clk_period;
		Addr <=  "0001110101000";
		Trees_din <= x"5bfef604";
		wait for Clk_period;
		Addr <=  "0001110101001";
		Trees_din <= x"00510fc5";
		wait for Clk_period;
		Addr <=  "0001110101010";
		Trees_din <= x"ff540fc5";
		wait for Clk_period;
		Addr <=  "0001110101011";
		Trees_din <= x"9bffee08";
		wait for Clk_period;
		Addr <=  "0001110101100";
		Trees_din <= x"e8feb304";
		wait for Clk_period;
		Addr <=  "0001110101101";
		Trees_din <= x"00a90fc5";
		wait for Clk_period;
		Addr <=  "0001110101110";
		Trees_din <= x"ff9a0fc5";
		wait for Clk_period;
		Addr <=  "0001110101111";
		Trees_din <= x"eaff6104";
		wait for Clk_period;
		Addr <=  "0001110110000";
		Trees_din <= x"ffec0fc5";
		wait for Clk_period;
		Addr <=  "0001110110001";
		Trees_din <= x"01330fc5";
		wait for Clk_period;
		Addr <=  "0001110110010";
		Trees_din <= x"7efebc40";
		wait for Clk_period;
		Addr <=  "0001110110011";
		Trees_din <= x"00ffce20";
		wait for Clk_period;
		Addr <=  "0001110110100";
		Trees_din <= x"c8000310";
		wait for Clk_period;
		Addr <=  "0001110110101";
		Trees_din <= x"96fef808";
		wait for Clk_period;
		Addr <=  "0001110110110";
		Trees_din <= x"86ffcb04";
		wait for Clk_period;
		Addr <=  "0001110110111";
		Trees_din <= x"00c40fc5";
		wait for Clk_period;
		Addr <=  "0001110111000";
		Trees_din <= x"ff720fc5";
		wait for Clk_period;
		Addr <=  "0001110111001";
		Trees_din <= x"6e004204";
		wait for Clk_period;
		Addr <=  "0001110111010";
		Trees_din <= x"ffee0fc5";
		wait for Clk_period;
		Addr <=  "0001110111011";
		Trees_din <= x"00550fc5";
		wait for Clk_period;
		Addr <=  "0001110111100";
		Trees_din <= x"80ffbb08";
		wait for Clk_period;
		Addr <=  "0001110111101";
		Trees_din <= x"82ff2a04";
		wait for Clk_period;
		Addr <=  "0001110111110";
		Trees_din <= x"00570fc5";
		wait for Clk_period;
		Addr <=  "0001110111111";
		Trees_din <= x"00b60fc5";
		wait for Clk_period;
		Addr <=  "0001111000000";
		Trees_din <= x"5a006404";
		wait for Clk_period;
		Addr <=  "0001111000001";
		Trees_din <= x"007e0fc5";
		wait for Clk_period;
		Addr <=  "0001111000010";
		Trees_din <= x"ffd30fc5";
		wait for Clk_period;
		Addr <=  "0001111000011";
		Trees_din <= x"cafe7010";
		wait for Clk_period;
		Addr <=  "0001111000100";
		Trees_din <= x"eaff6d08";
		wait for Clk_period;
		Addr <=  "0001111000101";
		Trees_din <= x"5bff9f04";
		wait for Clk_period;
		Addr <=  "0001111000110";
		Trees_din <= x"00ad0fc5";
		wait for Clk_period;
		Addr <=  "0001111000111";
		Trees_din <= x"ffb00fc5";
		wait for Clk_period;
		Addr <=  "0001111001000";
		Trees_din <= x"0affd904";
		wait for Clk_period;
		Addr <=  "0001111001001";
		Trees_din <= x"00a40fc5";
		wait for Clk_period;
		Addr <=  "0001111001010";
		Trees_din <= x"ffc10fc5";
		wait for Clk_period;
		Addr <=  "0001111001011";
		Trees_din <= x"d600fb08";
		wait for Clk_period;
		Addr <=  "0001111001100";
		Trees_din <= x"38003a04";
		wait for Clk_period;
		Addr <=  "0001111001101";
		Trees_din <= x"ff5d0fc5";
		wait for Clk_period;
		Addr <=  "0001111001110";
		Trees_din <= x"003e0fc5";
		wait for Clk_period;
		Addr <=  "0001111001111";
		Trees_din <= x"07011904";
		wait for Clk_period;
		Addr <=  "0001111010000";
		Trees_din <= x"ffcd0fc5";
		wait for Clk_period;
		Addr <=  "0001111010001";
		Trees_din <= x"00930fc5";
		wait for Clk_period;
		Addr <=  "0001111010010";
		Trees_din <= x"3bff9320";
		wait for Clk_period;
		Addr <=  "0001111010011";
		Trees_din <= x"71000710";
		wait for Clk_period;
		Addr <=  "0001111010100";
		Trees_din <= x"36ff9a08";
		wait for Clk_period;
		Addr <=  "0001111010101";
		Trees_din <= x"8c00c004";
		wait for Clk_period;
		Addr <=  "0001111010110";
		Trees_din <= x"ffc90fc5";
		wait for Clk_period;
		Addr <=  "0001111010111";
		Trees_din <= x"00870fc5";
		wait for Clk_period;
		Addr <=  "0001111011000";
		Trees_din <= x"6fffc304";
		wait for Clk_period;
		Addr <=  "0001111011001";
		Trees_din <= x"00040fc5";
		wait for Clk_period;
		Addr <=  "0001111011010";
		Trees_din <= x"00950fc5";
		wait for Clk_period;
		Addr <=  "0001111011011";
		Trees_din <= x"22ffb208";
		wait for Clk_period;
		Addr <=  "0001111011100";
		Trees_din <= x"d700e204";
		wait for Clk_period;
		Addr <=  "0001111011101";
		Trees_din <= x"ffa20fc5";
		wait for Clk_period;
		Addr <=  "0001111011110";
		Trees_din <= x"00b10fc5";
		wait for Clk_period;
		Addr <=  "0001111011111";
		Trees_din <= x"24fffd04";
		wait for Clk_period;
		Addr <=  "0001111100000";
		Trees_din <= x"01250fc5";
		wait for Clk_period;
		Addr <=  "0001111100001";
		Trees_din <= x"ff970fc5";
		wait for Clk_period;
		Addr <=  "0001111100010";
		Trees_din <= x"ee000110";
		wait for Clk_period;
		Addr <=  "0001111100011";
		Trees_din <= x"12ff6608";
		wait for Clk_period;
		Addr <=  "0001111100100";
		Trees_din <= x"19ff3204";
		wait for Clk_period;
		Addr <=  "0001111100101";
		Trees_din <= x"008e0fc5";
		wait for Clk_period;
		Addr <=  "0001111100110";
		Trees_din <= x"ff830fc5";
		wait for Clk_period;
		Addr <=  "0001111100111";
		Trees_din <= x"34ffe104";
		wait for Clk_period;
		Addr <=  "0001111101000";
		Trees_din <= x"fffc0fc5";
		wait for Clk_period;
		Addr <=  "0001111101001";
		Trees_din <= x"00cb0fc5";
		wait for Clk_period;
		Addr <=  "0001111101010";
		Trees_din <= x"0a001b08";
		wait for Clk_period;
		Addr <=  "0001111101011";
		Trees_din <= x"b4febf04";
		wait for Clk_period;
		Addr <=  "0001111101100";
		Trees_din <= x"ffaa0fc5";
		wait for Clk_period;
		Addr <=  "0001111101101";
		Trees_din <= x"008e0fc5";
		wait for Clk_period;
		Addr <=  "0001111101110";
		Trees_din <= x"0a00b504";
		wait for Clk_period;
		Addr <=  "0001111101111";
		Trees_din <= x"ff520fc5";
		wait for Clk_period;
		Addr <=  "0001111110000";
		Trees_din <= x"00490fc5";
		wait for Clk_period;
		Addr <=  "0001111110001";
		Trees_din <= x"36fee958";
		wait for Clk_period;
		Addr <=  "0001111110010";
		Trees_din <= x"70feea2c";
		wait for Clk_period;
		Addr <=  "0001111110011";
		Trees_din <= x"dfff3314";
		wait for Clk_period;
		Addr <=  "0001111110100";
		Trees_din <= x"18ff110c";
		wait for Clk_period;
		Addr <=  "0001111110101";
		Trees_din <= x"9aff5b04";
		wait for Clk_period;
		Addr <=  "0001111110110";
		Trees_din <= x"ff751159";
		wait for Clk_period;
		Addr <=  "0001111110111";
		Trees_din <= x"75005604";
		wait for Clk_period;
		Addr <=  "0001111111000";
		Trees_din <= x"00c41159";
		wait for Clk_period;
		Addr <=  "0001111111001";
		Trees_din <= x"002c1159";
		wait for Clk_period;
		Addr <=  "0001111111010";
		Trees_din <= x"28fe5104";
		wait for Clk_period;
		Addr <=  "0001111111011";
		Trees_din <= x"002f1159";
		wait for Clk_period;
		Addr <=  "0001111111100";
		Trees_din <= x"ff5b1159";
		wait for Clk_period;
		Addr <=  "0001111111101";
		Trees_din <= x"b2003c10";
		wait for Clk_period;
		Addr <=  "0001111111110";
		Trees_din <= x"0fff8608";
		wait for Clk_period;
		Addr <=  "0001111111111";
		Trees_din <= x"09ffea04";
		wait for Clk_period;
		Addr <=  "0010000000000";
		Trees_din <= x"ff8c1159";
		wait for Clk_period;
		Addr <=  "0010000000001";
		Trees_din <= x"006d1159";
		wait for Clk_period;
		Addr <=  "0010000000010";
		Trees_din <= x"f5003b04";
		wait for Clk_period;
		Addr <=  "0010000000011";
		Trees_din <= x"00c71159";
		wait for Clk_period;
		Addr <=  "0010000000100";
		Trees_din <= x"ffe11159";
		wait for Clk_period;
		Addr <=  "0010000000101";
		Trees_din <= x"56ff5f04";
		wait for Clk_period;
		Addr <=  "0010000000110";
		Trees_din <= x"000f1159";
		wait for Clk_period;
		Addr <=  "0010000000111";
		Trees_din <= x"ff601159";
		wait for Clk_period;
		Addr <=  "0010000001000";
		Trees_din <= x"18011020";
		wait for Clk_period;
		Addr <=  "0010000001001";
		Trees_din <= x"1f003210";
		wait for Clk_period;
		Addr <=  "0010000001010";
		Trees_din <= x"effec408";
		wait for Clk_period;
		Addr <=  "0010000001011";
		Trees_din <= x"a4ffa104";
		wait for Clk_period;
		Addr <=  "0010000001100";
		Trees_din <= x"ff851159";
		wait for Clk_period;
		Addr <=  "0010000001101";
		Trees_din <= x"00b51159";
		wait for Clk_period;
		Addr <=  "0010000001110";
		Trees_din <= x"44ff0f04";
		wait for Clk_period;
		Addr <=  "0010000001111";
		Trees_din <= x"00241159";
		wait for Clk_period;
		Addr <=  "0010000010000";
		Trees_din <= x"ff591159";
		wait for Clk_period;
		Addr <=  "0010000010001";
		Trees_din <= x"6d003908";
		wait for Clk_period;
		Addr <=  "0010000010010";
		Trees_din <= x"33fef104";
		wait for Clk_period;
		Addr <=  "0010000010011";
		Trees_din <= x"006b1159";
		wait for Clk_period;
		Addr <=  "0010000010100";
		Trees_din <= x"ff761159";
		wait for Clk_period;
		Addr <=  "0010000010101";
		Trees_din <= x"9bff5104";
		wait for Clk_period;
		Addr <=  "0010000010110";
		Trees_din <= x"00d81159";
		wait for Clk_period;
		Addr <=  "0010000010111";
		Trees_din <= x"ff9c1159";
		wait for Clk_period;
		Addr <=  "0010000011000";
		Trees_din <= x"c1fef708";
		wait for Clk_period;
		Addr <=  "0010000011001";
		Trees_din <= x"ac000104";
		wait for Clk_period;
		Addr <=  "0010000011010";
		Trees_din <= x"00a31159";
		wait for Clk_period;
		Addr <=  "0010000011011";
		Trees_din <= x"ff601159";
		wait for Clk_period;
		Addr <=  "0010000011100";
		Trees_din <= x"00e11159";
		wait for Clk_period;
		Addr <=  "0010000011101";
		Trees_din <= x"3d000034";
		wait for Clk_period;
		Addr <=  "0010000011110";
		Trees_din <= x"32ffb720";
		wait for Clk_period;
		Addr <=  "0010000011111";
		Trees_din <= x"9fff7810";
		wait for Clk_period;
		Addr <=  "0010000100000";
		Trees_din <= x"0d001c08";
		wait for Clk_period;
		Addr <=  "0010000100001";
		Trees_din <= x"f5007a04";
		wait for Clk_period;
		Addr <=  "0010000100010";
		Trees_din <= x"00651159";
		wait for Clk_period;
		Addr <=  "0010000100011";
		Trees_din <= x"ffd71159";
		wait for Clk_period;
		Addr <=  "0010000100100";
		Trees_din <= x"36ff3a04";
		wait for Clk_period;
		Addr <=  "0010000100101";
		Trees_din <= x"008d1159";
		wait for Clk_period;
		Addr <=  "0010000100110";
		Trees_din <= x"ffab1159";
		wait for Clk_period;
		Addr <=  "0010000100111";
		Trees_din <= x"25007008";
		wait for Clk_period;
		Addr <=  "0010000101000";
		Trees_din <= x"cafdaa04";
		wait for Clk_period;
		Addr <=  "0010000101001";
		Trees_din <= x"009e1159";
		wait for Clk_period;
		Addr <=  "0010000101010";
		Trees_din <= x"fff01159";
		wait for Clk_period;
		Addr <=  "0010000101011";
		Trees_din <= x"51008e04";
		wait for Clk_period;
		Addr <=  "0010000101100";
		Trees_din <= x"00811159";
		wait for Clk_period;
		Addr <=  "0010000101101";
		Trees_din <= x"ff851159";
		wait for Clk_period;
		Addr <=  "0010000101110";
		Trees_din <= x"0700960c";
		wait for Clk_period;
		Addr <=  "0010000101111";
		Trees_din <= x"cc004708";
		wait for Clk_period;
		Addr <=  "0010000110000";
		Trees_din <= x"48ff7e04";
		wait for Clk_period;
		Addr <=  "0010000110001";
		Trees_din <= x"003c1159";
		wait for Clk_period;
		Addr <=  "0010000110010";
		Trees_din <= x"ff6e1159";
		wait for Clk_period;
		Addr <=  "0010000110011";
		Trees_din <= x"00a11159";
		wait for Clk_period;
		Addr <=  "0010000110100";
		Trees_din <= x"d0007404";
		wait for Clk_period;
		Addr <=  "0010000110101";
		Trees_din <= x"fff11159";
		wait for Clk_period;
		Addr <=  "0010000110110";
		Trees_din <= x"00e61159";
		wait for Clk_period;
		Addr <=  "0010000110111";
		Trees_din <= x"7affa420";
		wait for Clk_period;
		Addr <=  "0010000111000";
		Trees_din <= x"85ff9f10";
		wait for Clk_period;
		Addr <=  "0010000111001";
		Trees_din <= x"72002f08";
		wait for Clk_period;
		Addr <=  "0010000111010";
		Trees_din <= x"0900b504";
		wait for Clk_period;
		Addr <=  "0010000111011";
		Trees_din <= x"ffda1159";
		wait for Clk_period;
		Addr <=  "0010000111100";
		Trees_din <= x"00f21159";
		wait for Clk_period;
		Addr <=  "0010000111101";
		Trees_din <= x"6e004204";
		wait for Clk_period;
		Addr <=  "0010000111110";
		Trees_din <= x"ffe31159";
		wait for Clk_period;
		Addr <=  "0010000111111";
		Trees_din <= x"00ab1159";
		wait for Clk_period;
		Addr <=  "0010001000000";
		Trees_din <= x"19feae08";
		wait for Clk_period;
		Addr <=  "0010001000001";
		Trees_din <= x"85ffe404";
		wait for Clk_period;
		Addr <=  "0010001000010";
		Trees_din <= x"010c1159";
		wait for Clk_period;
		Addr <=  "0010001000011";
		Trees_din <= x"ff9f1159";
		wait for Clk_period;
		Addr <=  "0010001000100";
		Trees_din <= x"40009f04";
		wait for Clk_period;
		Addr <=  "0010001000101";
		Trees_din <= x"ff901159";
		wait for Clk_period;
		Addr <=  "0010001000110";
		Trees_din <= x"008e1159";
		wait for Clk_period;
		Addr <=  "0010001000111";
		Trees_din <= x"5dff8c10";
		wait for Clk_period;
		Addr <=  "0010001001000";
		Trees_din <= x"c5ff7108";
		wait for Clk_period;
		Addr <=  "0010001001001";
		Trees_din <= x"83ff1204";
		wait for Clk_period;
		Addr <=  "0010001001010";
		Trees_din <= x"003c1159";
		wait for Clk_period;
		Addr <=  "0010001001011";
		Trees_din <= x"00e01159";
		wait for Clk_period;
		Addr <=  "0010001001100";
		Trees_din <= x"87ff5a04";
		wait for Clk_period;
		Addr <=  "0010001001101";
		Trees_din <= x"00641159";
		wait for Clk_period;
		Addr <=  "0010001001110";
		Trees_din <= x"ff621159";
		wait for Clk_period;
		Addr <=  "0010001001111";
		Trees_din <= x"d8004308";
		wait for Clk_period;
		Addr <=  "0010001010000";
		Trees_din <= x"76000504";
		wait for Clk_period;
		Addr <=  "0010001010001";
		Trees_din <= x"ffc41159";
		wait for Clk_period;
		Addr <=  "0010001010010";
		Trees_din <= x"00521159";
		wait for Clk_period;
		Addr <=  "0010001010011";
		Trees_din <= x"30ffe304";
		wait for Clk_period;
		Addr <=  "0010001010100";
		Trees_din <= x"00801159";
		wait for Clk_period;
		Addr <=  "0010001010101";
		Trees_din <= x"ffea1159";
		wait for Clk_period;
		Addr <=  "0010001010110";
		Trees_din <= x"cf001364";
		wait for Clk_period;
		Addr <=  "0010001010111";
		Trees_din <= x"95fec328";
		wait for Clk_period;
		Addr <=  "0010001011000";
		Trees_din <= x"a0ff4614";
		wait for Clk_period;
		Addr <=  "0010001011001";
		Trees_din <= x"cbff0604";
		wait for Clk_period;
		Addr <=  "0010001011010";
		Trees_din <= x"ff6c12fd";
		wait for Clk_period;
		Addr <=  "0010001011011";
		Trees_din <= x"36ff5c08";
		wait for Clk_period;
		Addr <=  "0010001011100";
		Trees_din <= x"6e008604";
		wait for Clk_period;
		Addr <=  "0010001011101";
		Trees_din <= x"ffdb12fd";
		wait for Clk_period;
		Addr <=  "0010001011110";
		Trees_din <= x"008312fd";
		wait for Clk_period;
		Addr <=  "0010001011111";
		Trees_din <= x"66ff6604";
		wait for Clk_period;
		Addr <=  "0010001100000";
		Trees_din <= x"ffc312fd";
		wait for Clk_period;
		Addr <=  "0010001100001";
		Trees_din <= x"00bf12fd";
		wait for Clk_period;
		Addr <=  "0010001100010";
		Trees_din <= x"8dfe0a04";
		wait for Clk_period;
		Addr <=  "0010001100011";
		Trees_din <= x"007f12fd";
		wait for Clk_period;
		Addr <=  "0010001100100";
		Trees_din <= x"6d00b408";
		wait for Clk_period;
		Addr <=  "0010001100101";
		Trees_din <= x"25ff9f04";
		wait for Clk_period;
		Addr <=  "0010001100110";
		Trees_din <= x"ffd512fd";
		wait for Clk_period;
		Addr <=  "0010001100111";
		Trees_din <= x"ff5312fd";
		wait for Clk_period;
		Addr <=  "0010001101000";
		Trees_din <= x"f0ffa404";
		wait for Clk_period;
		Addr <=  "0010001101001";
		Trees_din <= x"fff912fd";
		wait for Clk_period;
		Addr <=  "0010001101010";
		Trees_din <= x"008312fd";
		wait for Clk_period;
		Addr <=  "0010001101011";
		Trees_din <= x"4000021c";
		wait for Clk_period;
		Addr <=  "0010001101100";
		Trees_din <= x"61ff6c0c";
		wait for Clk_period;
		Addr <=  "0010001101101";
		Trees_din <= x"6dff9d04";
		wait for Clk_period;
		Addr <=  "0010001101110";
		Trees_din <= x"004b12fd";
		wait for Clk_period;
		Addr <=  "0010001101111";
		Trees_din <= x"03008c04";
		wait for Clk_period;
		Addr <=  "0010001110000";
		Trees_din <= x"ff5612fd";
		wait for Clk_period;
		Addr <=  "0010001110001";
		Trees_din <= x"fff912fd";
		wait for Clk_period;
		Addr <=  "0010001110010";
		Trees_din <= x"6a000408";
		wait for Clk_period;
		Addr <=  "0010001110011";
		Trees_din <= x"0fff6f04";
		wait for Clk_period;
		Addr <=  "0010001110100";
		Trees_din <= x"ff7412fd";
		wait for Clk_period;
		Addr <=  "0010001110101";
		Trees_din <= x"000812fd";
		wait for Clk_period;
		Addr <=  "0010001110110";
		Trees_din <= x"69ff2504";
		wait for Clk_period;
		Addr <=  "0010001110111";
		Trees_din <= x"ff8912fd";
		wait for Clk_period;
		Addr <=  "0010001111000";
		Trees_din <= x"00f712fd";
		wait for Clk_period;
		Addr <=  "0010001111001";
		Trees_din <= x"5bff9310";
		wait for Clk_period;
		Addr <=  "0010001111010";
		Trees_din <= x"34ffe508";
		wait for Clk_period;
		Addr <=  "0010001111011";
		Trees_din <= x"d500b704";
		wait for Clk_period;
		Addr <=  "0010001111100";
		Trees_din <= x"ffb212fd";
		wait for Clk_period;
		Addr <=  "0010001111101";
		Trees_din <= x"007b12fd";
		wait for Clk_period;
		Addr <=  "0010001111110";
		Trees_din <= x"84ffe604";
		wait for Clk_period;
		Addr <=  "0010001111111";
		Trees_din <= x"005712fd";
		wait for Clk_period;
		Addr <=  "0010010000000";
		Trees_din <= x"fff212fd";
		wait for Clk_period;
		Addr <=  "0010010000001";
		Trees_din <= x"bcfef008";
		wait for Clk_period;
		Addr <=  "0010010000010";
		Trees_din <= x"30001604";
		wait for Clk_period;
		Addr <=  "0010010000011";
		Trees_din <= x"002412fd";
		wait for Clk_period;
		Addr <=  "0010010000100";
		Trees_din <= x"ff8212fd";
		wait for Clk_period;
		Addr <=  "0010010000101";
		Trees_din <= x"09009a04";
		wait for Clk_period;
		Addr <=  "0010010000110";
		Trees_din <= x"ff7312fd";
		wait for Clk_period;
		Addr <=  "0010010000111";
		Trees_din <= x"007c12fd";
		wait for Clk_period;
		Addr <=  "0010010001000";
		Trees_din <= x"a1ffab3c";
		wait for Clk_period;
		Addr <=  "0010010001001";
		Trees_din <= x"61ffe220";
		wait for Clk_period;
		Addr <=  "0010010001010";
		Trees_din <= x"1dff0b10";
		wait for Clk_period;
		Addr <=  "0010010001011";
		Trees_din <= x"17ffe608";
		wait for Clk_period;
		Addr <=  "0010010001100";
		Trees_din <= x"81ffd104";
		wait for Clk_period;
		Addr <=  "0010010001101";
		Trees_din <= x"006812fd";
		wait for Clk_period;
		Addr <=  "0010010001110";
		Trees_din <= x"fff012fd";
		wait for Clk_period;
		Addr <=  "0010010001111";
		Trees_din <= x"d2ff8404";
		wait for Clk_period;
		Addr <=  "0010010010000";
		Trees_din <= x"ffe912fd";
		wait for Clk_period;
		Addr <=  "0010010010001";
		Trees_din <= x"00f812fd";
		wait for Clk_period;
		Addr <=  "0010010010010";
		Trees_din <= x"d3fe6208";
		wait for Clk_period;
		Addr <=  "0010010010011";
		Trees_din <= x"0500bc04";
		wait for Clk_period;
		Addr <=  "0010010010100";
		Trees_din <= x"ff8012fd";
		wait for Clk_period;
		Addr <=  "0010010010101";
		Trees_din <= x"007612fd";
		wait for Clk_period;
		Addr <=  "0010010010110";
		Trees_din <= x"31ff6404";
		wait for Clk_period;
		Addr <=  "0010010010111";
		Trees_din <= x"fffc12fd";
		wait for Clk_period;
		Addr <=  "0010010011000";
		Trees_din <= x"005c12fd";
		wait for Clk_period;
		Addr <=  "0010010011001";
		Trees_din <= x"74004d10";
		wait for Clk_period;
		Addr <=  "0010010011010";
		Trees_din <= x"71ff1f08";
		wait for Clk_period;
		Addr <=  "0010010011011";
		Trees_din <= x"1eff7204";
		wait for Clk_period;
		Addr <=  "0010010011100";
		Trees_din <= x"009f12fd";
		wait for Clk_period;
		Addr <=  "0010010011101";
		Trees_din <= x"001812fd";
		wait for Clk_period;
		Addr <=  "0010010011110";
		Trees_din <= x"c3ffbf04";
		wait for Clk_period;
		Addr <=  "0010010011111";
		Trees_din <= x"003012fd";
		wait for Clk_period;
		Addr <=  "0010010100000";
		Trees_din <= x"00be12fd";
		wait for Clk_period;
		Addr <=  "0010010100001";
		Trees_din <= x"e2ff7608";
		wait for Clk_period;
		Addr <=  "0010010100010";
		Trees_din <= x"29ffbe04";
		wait for Clk_period;
		Addr <=  "0010010100011";
		Trees_din <= x"ff5912fd";
		wait for Clk_period;
		Addr <=  "0010010100100";
		Trees_din <= x"ffe012fd";
		wait for Clk_period;
		Addr <=  "0010010100101";
		Trees_din <= x"007a12fd";
		wait for Clk_period;
		Addr <=  "0010010100110";
		Trees_din <= x"2bff3914";
		wait for Clk_period;
		Addr <=  "0010010100111";
		Trees_din <= x"f0ff900c";
		wait for Clk_period;
		Addr <=  "0010010101000";
		Trees_din <= x"4effeb08";
		wait for Clk_period;
		Addr <=  "0010010101001";
		Trees_din <= x"1e003304";
		wait for Clk_period;
		Addr <=  "0010010101010";
		Trees_din <= x"010912fd";
		wait for Clk_period;
		Addr <=  "0010010101011";
		Trees_din <= x"fff812fd";
		wait for Clk_period;
		Addr <=  "0010010101100";
		Trees_din <= x"ffd912fd";
		wait for Clk_period;
		Addr <=  "0010010101101";
		Trees_din <= x"a0feaa04";
		wait for Clk_period;
		Addr <=  "0010010101110";
		Trees_din <= x"003512fd";
		wait for Clk_period;
		Addr <=  "0010010101111";
		Trees_din <= x"ff8412fd";
		wait for Clk_period;
		Addr <=  "0010010110000";
		Trees_din <= x"42ff2710";
		wait for Clk_period;
		Addr <=  "0010010110001";
		Trees_din <= x"1bff8508";
		wait for Clk_period;
		Addr <=  "0010010110010";
		Trees_din <= x"8bffec04";
		wait for Clk_period;
		Addr <=  "0010010110011";
		Trees_din <= x"000c12fd";
		wait for Clk_period;
		Addr <=  "0010010110100";
		Trees_din <= x"ff7712fd";
		wait for Clk_period;
		Addr <=  "0010010110101";
		Trees_din <= x"70ff5704";
		wait for Clk_period;
		Addr <=  "0010010110110";
		Trees_din <= x"00bf12fd";
		wait for Clk_period;
		Addr <=  "0010010110111";
		Trees_din <= x"ff8f12fd";
		wait for Clk_period;
		Addr <=  "0010010111000";
		Trees_din <= x"a6feee08";
		wait for Clk_period;
		Addr <=  "0010010111001";
		Trees_din <= x"70ff0104";
		wait for Clk_period;
		Addr <=  "0010010111010";
		Trees_din <= x"00b212fd";
		wait for Clk_period;
		Addr <=  "0010010111011";
		Trees_din <= x"ff9b12fd";
		wait for Clk_period;
		Addr <=  "0010010111100";
		Trees_din <= x"41ffa304";
		wait for Clk_period;
		Addr <=  "0010010111101";
		Trees_din <= x"ff7a12fd";
		wait for Clk_period;
		Addr <=  "0010010111110";
		Trees_din <= x"005212fd";
		wait for Clk_period;
		Addr <=  "0010010111111";
		Trees_din <= x"6f003e60";
		wait for Clk_period;
		Addr <=  "0010011000000";
		Trees_din <= x"6d007040";
		wait for Clk_period;
		Addr <=  "0010011000001";
		Trees_din <= x"72005220";
		wait for Clk_period;
		Addr <=  "0010011000010";
		Trees_din <= x"1efee610";
		wait for Clk_period;
		Addr <=  "0010011000011";
		Trees_din <= x"60ffa408";
		wait for Clk_period;
		Addr <=  "0010011000100";
		Trees_din <= x"f6ff0f04";
		wait for Clk_period;
		Addr <=  "0010011000101";
		Trees_din <= x"005d1409";
		wait for Clk_period;
		Addr <=  "0010011000110";
		Trees_din <= x"ff681409";
		wait for Clk_period;
		Addr <=  "0010011000111";
		Trees_din <= x"b4ff6b04";
		wait for Clk_period;
		Addr <=  "0010011001000";
		Trees_din <= x"00de1409";
		wait for Clk_period;
		Addr <=  "0010011001001";
		Trees_din <= x"fff71409";
		wait for Clk_period;
		Addr <=  "0010011001010";
		Trees_din <= x"64ff6608";
		wait for Clk_period;
		Addr <=  "0010011001011";
		Trees_din <= x"34fff804";
		wait for Clk_period;
		Addr <=  "0010011001100";
		Trees_din <= x"ffb91409";
		wait for Clk_period;
		Addr <=  "0010011001101";
		Trees_din <= x"fff81409";
		wait for Clk_period;
		Addr <=  "0010011001110";
		Trees_din <= x"f3ff0404";
		wait for Clk_period;
		Addr <=  "0010011001111";
		Trees_din <= x"00341409";
		wait for Clk_period;
		Addr <=  "0010011010000";
		Trees_din <= x"ffdd1409";
		wait for Clk_period;
		Addr <=  "0010011010001";
		Trees_din <= x"87ff2f10";
		wait for Clk_period;
		Addr <=  "0010011010010";
		Trees_din <= x"90fff508";
		wait for Clk_period;
		Addr <=  "0010011010011";
		Trees_din <= x"2dff3704";
		wait for Clk_period;
		Addr <=  "0010011010100";
		Trees_din <= x"00a11409";
		wait for Clk_period;
		Addr <=  "0010011010101";
		Trees_din <= x"fffc1409";
		wait for Clk_period;
		Addr <=  "0010011010110";
		Trees_din <= x"0400cb04";
		wait for Clk_period;
		Addr <=  "0010011010111";
		Trees_din <= x"ff6c1409";
		wait for Clk_period;
		Addr <=  "0010011011000";
		Trees_din <= x"00541409";
		wait for Clk_period;
		Addr <=  "0010011011001";
		Trees_din <= x"ebff4908";
		wait for Clk_period;
		Addr <=  "0010011011010";
		Trees_din <= x"c3001e04";
		wait for Clk_period;
		Addr <=  "0010011011011";
		Trees_din <= x"00051409";
		wait for Clk_period;
		Addr <=  "0010011011100";
		Trees_din <= x"00641409";
		wait for Clk_period;
		Addr <=  "0010011011101";
		Trees_din <= x"1b002704";
		wait for Clk_period;
		Addr <=  "0010011011110";
		Trees_din <= x"ff571409";
		wait for Clk_period;
		Addr <=  "0010011011111";
		Trees_din <= x"002d1409";
		wait for Clk_period;
		Addr <=  "0010011100000";
		Trees_din <= x"3d007614";
		wait for Clk_period;
		Addr <=  "0010011100001";
		Trees_din <= x"50fe2b04";
		wait for Clk_period;
		Addr <=  "0010011100010";
		Trees_din <= x"ff681409";
		wait for Clk_period;
		Addr <=  "0010011100011";
		Trees_din <= x"20ff4708";
		wait for Clk_period;
		Addr <=  "0010011100100";
		Trees_din <= x"7d000d04";
		wait for Clk_period;
		Addr <=  "0010011100101";
		Trees_din <= x"ffc61409";
		wait for Clk_period;
		Addr <=  "0010011100110";
		Trees_din <= x"00651409";
		wait for Clk_period;
		Addr <=  "0010011100111";
		Trees_din <= x"a0ff5e04";
		wait for Clk_period;
		Addr <=  "0010011101000";
		Trees_din <= x"00721409";
		wait for Clk_period;
		Addr <=  "0010011101001";
		Trees_din <= x"00031409";
		wait for Clk_period;
		Addr <=  "0010011101010";
		Trees_din <= x"5400cc08";
		wait for Clk_period;
		Addr <=  "0010011101011";
		Trees_din <= x"59ffe904";
		wait for Clk_period;
		Addr <=  "0010011101100";
		Trees_din <= x"ff601409";
		wait for Clk_period;
		Addr <=  "0010011101101";
		Trees_din <= x"00261409";
		wait for Clk_period;
		Addr <=  "0010011101110";
		Trees_din <= x"00811409";
		wait for Clk_period;
		Addr <=  "0010011101111";
		Trees_din <= x"f203b024";
		wait for Clk_period;
		Addr <=  "0010011110000";
		Trees_din <= x"05fffe10";
		wait for Clk_period;
		Addr <=  "0010011110001";
		Trees_din <= x"d3fef208";
		wait for Clk_period;
		Addr <=  "0010011110010";
		Trees_din <= x"d9ffcf04";
		wait for Clk_period;
		Addr <=  "0010011110011";
		Trees_din <= x"00de1409";
		wait for Clk_period;
		Addr <=  "0010011110100";
		Trees_din <= x"ff9b1409";
		wait for Clk_period;
		Addr <=  "0010011110101";
		Trees_din <= x"6cff2604";
		wait for Clk_period;
		Addr <=  "0010011110110";
		Trees_din <= x"ffec1409";
		wait for Clk_period;
		Addr <=  "0010011110111";
		Trees_din <= x"ff761409";
		wait for Clk_period;
		Addr <=  "0010011111000";
		Trees_din <= x"38fee004";
		wait for Clk_period;
		Addr <=  "0010011111001";
		Trees_din <= x"ff981409";
		wait for Clk_period;
		Addr <=  "0010011111010";
		Trees_din <= x"ccff3908";
		wait for Clk_period;
		Addr <=  "0010011111011";
		Trees_din <= x"30ff7804";
		wait for Clk_period;
		Addr <=  "0010011111100";
		Trees_din <= x"008e1409";
		wait for Clk_period;
		Addr <=  "0010011111101";
		Trees_din <= x"ff7b1409";
		wait for Clk_period;
		Addr <=  "0010011111110";
		Trees_din <= x"75008604";
		wait for Clk_period;
		Addr <=  "0010011111111";
		Trees_din <= x"00d51409";
		wait for Clk_period;
		Addr <=  "0010100000000";
		Trees_din <= x"00151409";
		wait for Clk_period;
		Addr <=  "0010100000001";
		Trees_din <= x"ff741409";
		wait for Clk_period;
		Addr <=  "0010100000010";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0010100000011";
		Trees_din <= x"60ffbe78";
		wait for Clk_period;
		Addr <=  "0010100000100";
		Trees_din <= x"54002638";
		wait for Clk_period;
		Addr <=  "0010100000101";
		Trees_din <= x"4700291c";
		wait for Clk_period;
		Addr <=  "0010100000110";
		Trees_din <= x"d7ffc20c";
		wait for Clk_period;
		Addr <=  "0010100000111";
		Trees_din <= x"bd002708";
		wait for Clk_period;
		Addr <=  "0010100001000";
		Trees_din <= x"c6ff6304";
		wait for Clk_period;
		Addr <=  "0010100001001";
		Trees_din <= x"ffbf15c1";
		wait for Clk_period;
		Addr <=  "0010100001010";
		Trees_din <= x"010615c1";
		wait for Clk_period;
		Addr <=  "0010100001011";
		Trees_din <= x"ff8615c1";
		wait for Clk_period;
		Addr <=  "0010100001100";
		Trees_din <= x"25005208";
		wait for Clk_period;
		Addr <=  "0010100001101";
		Trees_din <= x"f1ff7104";
		wait for Clk_period;
		Addr <=  "0010100001110";
		Trees_din <= x"ffe115c1";
		wait for Clk_period;
		Addr <=  "0010100001111";
		Trees_din <= x"ff7815c1";
		wait for Clk_period;
		Addr <=  "0010100010000";
		Trees_din <= x"abffc704";
		wait for Clk_period;
		Addr <=  "0010100010001";
		Trees_din <= x"00a415c1";
		wait for Clk_period;
		Addr <=  "0010100010010";
		Trees_din <= x"ffcd15c1";
		wait for Clk_period;
		Addr <=  "0010100010011";
		Trees_din <= x"0bff280c";
		wait for Clk_period;
		Addr <=  "0010100010100";
		Trees_din <= x"a2ff7204";
		wait for Clk_period;
		Addr <=  "0010100010101";
		Trees_din <= x"ffa115c1";
		wait for Clk_period;
		Addr <=  "0010100010110";
		Trees_din <= x"c8ffd704";
		wait for Clk_period;
		Addr <=  "0010100010111";
		Trees_din <= x"fff215c1";
		wait for Clk_period;
		Addr <=  "0010100011000";
		Trees_din <= x"011615c1";
		wait for Clk_period;
		Addr <=  "0010100011001";
		Trees_din <= x"5c000708";
		wait for Clk_period;
		Addr <=  "0010100011010";
		Trees_din <= x"64ff0f04";
		wait for Clk_period;
		Addr <=  "0010100011011";
		Trees_din <= x"ff7f15c1";
		wait for Clk_period;
		Addr <=  "0010100011100";
		Trees_din <= x"000415c1";
		wait for Clk_period;
		Addr <=  "0010100011101";
		Trees_din <= x"78ff6004";
		wait for Clk_period;
		Addr <=  "0010100011110";
		Trees_din <= x"009e15c1";
		wait for Clk_period;
		Addr <=  "0010100011111";
		Trees_din <= x"fff715c1";
		wait for Clk_period;
		Addr <=  "0010100100000";
		Trees_din <= x"24ff8f20";
		wait for Clk_period;
		Addr <=  "0010100100001";
		Trees_din <= x"89003c10";
		wait for Clk_period;
		Addr <=  "0010100100010";
		Trees_din <= x"4eff0908";
		wait for Clk_period;
		Addr <=  "0010100100011";
		Trees_din <= x"54006b04";
		wait for Clk_period;
		Addr <=  "0010100100100";
		Trees_din <= x"00dc15c1";
		wait for Clk_period;
		Addr <=  "0010100100101";
		Trees_din <= x"005515c1";
		wait for Clk_period;
		Addr <=  "0010100100110";
		Trees_din <= x"40001404";
		wait for Clk_period;
		Addr <=  "0010100100111";
		Trees_din <= x"fffb15c1";
		wait for Clk_period;
		Addr <=  "0010100101000";
		Trees_din <= x"005a15c1";
		wait for Clk_period;
		Addr <=  "0010100101001";
		Trees_din <= x"7afff508";
		wait for Clk_period;
		Addr <=  "0010100101010";
		Trees_din <= x"78ff4604";
		wait for Clk_period;
		Addr <=  "0010100101011";
		Trees_din <= x"002a15c1";
		wait for Clk_period;
		Addr <=  "0010100101100";
		Trees_din <= x"ffa015c1";
		wait for Clk_period;
		Addr <=  "0010100101101";
		Trees_din <= x"6c003104";
		wait for Clk_period;
		Addr <=  "0010100101110";
		Trees_din <= x"008015c1";
		wait for Clk_period;
		Addr <=  "0010100101111";
		Trees_din <= x"ff7515c1";
		wait for Clk_period;
		Addr <=  "0010100110000";
		Trees_din <= x"95ff7610";
		wait for Clk_period;
		Addr <=  "0010100110001";
		Trees_din <= x"2dff1508";
		wait for Clk_period;
		Addr <=  "0010100110010";
		Trees_din <= x"3a000404";
		wait for Clk_period;
		Addr <=  "0010100110011";
		Trees_din <= x"ffeb15c1";
		wait for Clk_period;
		Addr <=  "0010100110100";
		Trees_din <= x"006215c1";
		wait for Clk_period;
		Addr <=  "0010100110101";
		Trees_din <= x"19ff3704";
		wait for Clk_period;
		Addr <=  "0010100110110";
		Trees_din <= x"007d15c1";
		wait for Clk_period;
		Addr <=  "0010100110111";
		Trees_din <= x"001415c1";
		wait for Clk_period;
		Addr <=  "0010100111000";
		Trees_din <= x"34002c08";
		wait for Clk_period;
		Addr <=  "0010100111001";
		Trees_din <= x"cb006204";
		wait for Clk_period;
		Addr <=  "0010100111010";
		Trees_din <= x"ff8b15c1";
		wait for Clk_period;
		Addr <=  "0010100111011";
		Trees_din <= x"007515c1";
		wait for Clk_period;
		Addr <=  "0010100111100";
		Trees_din <= x"91ff4004";
		wait for Clk_period;
		Addr <=  "0010100111101";
		Trees_din <= x"00c815c1";
		wait for Clk_period;
		Addr <=  "0010100111110";
		Trees_din <= x"ffd615c1";
		wait for Clk_period;
		Addr <=  "0010100111111";
		Trees_din <= x"05000124";
		wait for Clk_period;
		Addr <=  "0010101000000";
		Trees_din <= x"4800001c";
		wait for Clk_period;
		Addr <=  "0010101000001";
		Trees_din <= x"24ff9c0c";
		wait for Clk_period;
		Addr <=  "0010101000010";
		Trees_din <= x"feffbd08";
		wait for Clk_period;
		Addr <=  "0010101000011";
		Trees_din <= x"5cffeb04";
		wait for Clk_period;
		Addr <=  "0010101000100";
		Trees_din <= x"00f815c1";
		wait for Clk_period;
		Addr <=  "0010101000101";
		Trees_din <= x"fff615c1";
		wait for Clk_period;
		Addr <=  "0010101000110";
		Trees_din <= x"ff8415c1";
		wait for Clk_period;
		Addr <=  "0010101000111";
		Trees_din <= x"1bffe908";
		wait for Clk_period;
		Addr <=  "0010101001000";
		Trees_din <= x"37ff2a04";
		wait for Clk_period;
		Addr <=  "0010101001001";
		Trees_din <= x"004715c1";
		wait for Clk_period;
		Addr <=  "0010101001010";
		Trees_din <= x"ff6215c1";
		wait for Clk_period;
		Addr <=  "0010101001011";
		Trees_din <= x"b6ff5004";
		wait for Clk_period;
		Addr <=  "0010101001100";
		Trees_din <= x"009615c1";
		wait for Clk_period;
		Addr <=  "0010101001101";
		Trees_din <= x"ffa515c1";
		wait for Clk_period;
		Addr <=  "0010101001110";
		Trees_din <= x"0d003004";
		wait for Clk_period;
		Addr <=  "0010101001111";
		Trees_din <= x"ff5615c1";
		wait for Clk_period;
		Addr <=  "0010101010000";
		Trees_din <= x"001d15c1";
		wait for Clk_period;
		Addr <=  "0010101010001";
		Trees_din <= x"e8ff9420";
		wait for Clk_period;
		Addr <=  "0010101010010";
		Trees_din <= x"7aff2b10";
		wait for Clk_period;
		Addr <=  "0010101010011";
		Trees_din <= x"97ff3a08";
		wait for Clk_period;
		Addr <=  "0010101010100";
		Trees_din <= x"c0ffad04";
		wait for Clk_period;
		Addr <=  "0010101010101";
		Trees_din <= x"ff5f15c1";
		wait for Clk_period;
		Addr <=  "0010101010110";
		Trees_din <= x"001b15c1";
		wait for Clk_period;
		Addr <=  "0010101010111";
		Trees_din <= x"ec000204";
		wait for Clk_period;
		Addr <=  "0010101011000";
		Trees_din <= x"00ac15c1";
		wait for Clk_period;
		Addr <=  "0010101011001";
		Trees_din <= x"ff8515c1";
		wait for Clk_period;
		Addr <=  "0010101011010";
		Trees_din <= x"32fece08";
		wait for Clk_period;
		Addr <=  "0010101011011";
		Trees_din <= x"5bff6604";
		wait for Clk_period;
		Addr <=  "0010101011100";
		Trees_din <= x"008915c1";
		wait for Clk_period;
		Addr <=  "0010101011101";
		Trees_din <= x"000815c1";
		wait for Clk_period;
		Addr <=  "0010101011110";
		Trees_din <= x"f0fe4504";
		wait for Clk_period;
		Addr <=  "0010101011111";
		Trees_din <= x"ff7d15c1";
		wait for Clk_period;
		Addr <=  "0010101100000";
		Trees_din <= x"00c015c1";
		wait for Clk_period;
		Addr <=  "0010101100001";
		Trees_din <= x"86fefa10";
		wait for Clk_period;
		Addr <=  "0010101100010";
		Trees_din <= x"c5ff2308";
		wait for Clk_period;
		Addr <=  "0010101100011";
		Trees_din <= x"c0ff8104";
		wait for Clk_period;
		Addr <=  "0010101100100";
		Trees_din <= x"005215c1";
		wait for Clk_period;
		Addr <=  "0010101100101";
		Trees_din <= x"ff8615c1";
		wait for Clk_period;
		Addr <=  "0010101100110";
		Trees_din <= x"e0ff9204";
		wait for Clk_period;
		Addr <=  "0010101100111";
		Trees_din <= x"005615c1";
		wait for Clk_period;
		Addr <=  "0010101101000";
		Trees_din <= x"00f015c1";
		wait for Clk_period;
		Addr <=  "0010101101001";
		Trees_din <= x"3dff6608";
		wait for Clk_period;
		Addr <=  "0010101101010";
		Trees_din <= x"bd001704";
		wait for Clk_period;
		Addr <=  "0010101101011";
		Trees_din <= x"00b715c1";
		wait for Clk_period;
		Addr <=  "0010101101100";
		Trees_din <= x"ffbf15c1";
		wait for Clk_period;
		Addr <=  "0010101101101";
		Trees_din <= x"5a00be04";
		wait for Clk_period;
		Addr <=  "0010101101110";
		Trees_din <= x"ffba15c1";
		wait for Clk_period;
		Addr <=  "0010101101111";
		Trees_din <= x"004d15c1";
		wait for Clk_period;
		Addr <=  "0010101110000";
		Trees_din <= x"6f003e70";
		wait for Clk_period;
		Addr <=  "0010101110001";
		Trees_din <= x"a0ff6534";
		wait for Clk_period;
		Addr <=  "0010101110010";
		Trees_din <= x"1eff9914";
		wait for Clk_period;
		Addr <=  "0010101110011";
		Trees_din <= x"f5009d10";
		wait for Clk_period;
		Addr <=  "0010101110100";
		Trees_din <= x"8cfed008";
		wait for Clk_period;
		Addr <=  "0010101110101";
		Trees_din <= x"d1ff5704";
		wait for Clk_period;
		Addr <=  "0010101110110";
		Trees_din <= x"ff7416f5";
		wait for Clk_period;
		Addr <=  "0010101110111";
		Trees_din <= x"006816f5";
		wait for Clk_period;
		Addr <=  "0010101111000";
		Trees_din <= x"bcffc804";
		wait for Clk_period;
		Addr <=  "0010101111001";
		Trees_din <= x"003716f5";
		wait for Clk_period;
		Addr <=  "0010101111010";
		Trees_din <= x"ffba16f5";
		wait for Clk_period;
		Addr <=  "0010101111011";
		Trees_din <= x"ff6716f5";
		wait for Clk_period;
		Addr <=  "0010101111100";
		Trees_din <= x"74001010";
		wait for Clk_period;
		Addr <=  "0010101111101";
		Trees_din <= x"ebff5b08";
		wait for Clk_period;
		Addr <=  "0010101111110";
		Trees_din <= x"9bff3d04";
		wait for Clk_period;
		Addr <=  "0010101111111";
		Trees_din <= x"003b16f5";
		wait for Clk_period;
		Addr <=  "0010110000000";
		Trees_din <= x"ffff16f5";
		wait for Clk_period;
		Addr <=  "0010110000001";
		Trees_din <= x"6bfe5604";
		wait for Clk_period;
		Addr <=  "0010110000010";
		Trees_din <= x"006f16f5";
		wait for Clk_period;
		Addr <=  "0010110000011";
		Trees_din <= x"ff7416f5";
		wait for Clk_period;
		Addr <=  "0010110000100";
		Trees_din <= x"cafdaa08";
		wait for Clk_period;
		Addr <=  "0010110000101";
		Trees_din <= x"45ff1004";
		wait for Clk_period;
		Addr <=  "0010110000110";
		Trees_din <= x"00a516f5";
		wait for Clk_period;
		Addr <=  "0010110000111";
		Trees_din <= x"ffc016f5";
		wait for Clk_period;
		Addr <=  "0010110001000";
		Trees_din <= x"3affe404";
		wait for Clk_period;
		Addr <=  "0010110001001";
		Trees_din <= x"ffb716f5";
		wait for Clk_period;
		Addr <=  "0010110001010";
		Trees_din <= x"003116f5";
		wait for Clk_period;
		Addr <=  "0010110001011";
		Trees_din <= x"0fff941c";
		wait for Clk_period;
		Addr <=  "0010110001100";
		Trees_din <= x"93003d10";
		wait for Clk_period;
		Addr <=  "0010110001101";
		Trees_din <= x"d700cf08";
		wait for Clk_period;
		Addr <=  "0010110001110";
		Trees_din <= x"08011a04";
		wait for Clk_period;
		Addr <=  "0010110001111";
		Trees_din <= x"ff8316f5";
		wait for Clk_period;
		Addr <=  "0010110010000";
		Trees_din <= x"004d16f5";
		wait for Clk_period;
		Addr <=  "0010110010001";
		Trees_din <= x"97ff2d04";
		wait for Clk_period;
		Addr <=  "0010110010010";
		Trees_din <= x"ff9616f5";
		wait for Clk_period;
		Addr <=  "0010110010011";
		Trees_din <= x"008016f5";
		wait for Clk_period;
		Addr <=  "0010110010100";
		Trees_din <= x"eaffc808";
		wait for Clk_period;
		Addr <=  "0010110010101";
		Trees_din <= x"aeff5304";
		wait for Clk_period;
		Addr <=  "0010110010110";
		Trees_din <= x"00a616f5";
		wait for Clk_period;
		Addr <=  "0010110010111";
		Trees_din <= x"ffd316f5";
		wait for Clk_period;
		Addr <=  "0010110011000";
		Trees_din <= x"ff9c16f5";
		wait for Clk_period;
		Addr <=  "0010110011001";
		Trees_din <= x"09fff210";
		wait for Clk_period;
		Addr <=  "0010110011010";
		Trees_din <= x"1dff5008";
		wait for Clk_period;
		Addr <=  "0010110011011";
		Trees_din <= x"6fffec04";
		wait for Clk_period;
		Addr <=  "0010110011100";
		Trees_din <= x"ff7016f5";
		wait for Clk_period;
		Addr <=  "0010110011101";
		Trees_din <= x"003016f5";
		wait for Clk_period;
		Addr <=  "0010110011110";
		Trees_din <= x"08002104";
		wait for Clk_period;
		Addr <=  "0010110011111";
		Trees_din <= x"ff7a16f5";
		wait for Clk_period;
		Addr <=  "0010110100000";
		Trees_din <= x"006e16f5";
		wait for Clk_period;
		Addr <=  "0010110100001";
		Trees_din <= x"a8ff8108";
		wait for Clk_period;
		Addr <=  "0010110100010";
		Trees_din <= x"66000004";
		wait for Clk_period;
		Addr <=  "0010110100011";
		Trees_din <= x"ff9b16f5";
		wait for Clk_period;
		Addr <=  "0010110100100";
		Trees_din <= x"008b16f5";
		wait for Clk_period;
		Addr <=  "0010110100101";
		Trees_din <= x"25ffa804";
		wait for Clk_period;
		Addr <=  "0010110100110";
		Trees_din <= x"ffdb16f5";
		wait for Clk_period;
		Addr <=  "0010110100111";
		Trees_din <= x"00ce16f5";
		wait for Clk_period;
		Addr <=  "0010110101000";
		Trees_din <= x"8cff6710";
		wait for Clk_period;
		Addr <=  "0010110101001";
		Trees_din <= x"19ff6608";
		wait for Clk_period;
		Addr <=  "0010110101010";
		Trees_din <= x"ebfe8804";
		wait for Clk_period;
		Addr <=  "0010110101011";
		Trees_din <= x"002e16f5";
		wait for Clk_period;
		Addr <=  "0010110101100";
		Trees_din <= x"ff6316f5";
		wait for Clk_period;
		Addr <=  "0010110101101";
		Trees_din <= x"4dfe6004";
		wait for Clk_period;
		Addr <=  "0010110101110";
		Trees_din <= x"000016f5";
		wait for Clk_period;
		Addr <=  "0010110101111";
		Trees_din <= x"00c616f5";
		wait for Clk_period;
		Addr <=  "0010110110000";
		Trees_din <= x"38fef404";
		wait for Clk_period;
		Addr <=  "0010110110001";
		Trees_din <= x"ff9b16f5";
		wait for Clk_period;
		Addr <=  "0010110110010";
		Trees_din <= x"f6fe8e08";
		wait for Clk_period;
		Addr <=  "0010110110011";
		Trees_din <= x"38ff9a04";
		wait for Clk_period;
		Addr <=  "0010110110100";
		Trees_din <= x"ff8516f5";
		wait for Clk_period;
		Addr <=  "0010110110101";
		Trees_din <= x"004816f5";
		wait for Clk_period;
		Addr <=  "0010110110110";
		Trees_din <= x"baff0c08";
		wait for Clk_period;
		Addr <=  "0010110110111";
		Trees_din <= x"76ffaa04";
		wait for Clk_period;
		Addr <=  "0010110111000";
		Trees_din <= x"002f16f5";
		wait for Clk_period;
		Addr <=  "0010110111001";
		Trees_din <= x"ff9016f5";
		wait for Clk_period;
		Addr <=  "0010110111010";
		Trees_din <= x"04ffcc04";
		wait for Clk_period;
		Addr <=  "0010110111011";
		Trees_din <= x"ffa516f5";
		wait for Clk_period;
		Addr <=  "0010110111100";
		Trees_din <= x"00b916f5";
		wait for Clk_period;
		Addr <=  "0010110111101";
		Trees_din <= x"cf001574";
		wait for Clk_period;
		Addr <=  "0010110111110";
		Trees_din <= x"95fec338";
		wait for Clk_period;
		Addr <=  "0010110111111";
		Trees_din <= x"a0ff271c";
		wait for Clk_period;
		Addr <=  "0010111000000";
		Trees_din <= x"92ff0b0c";
		wait for Clk_period;
		Addr <=  "0010111000001";
		Trees_din <= x"f800c708";
		wait for Clk_period;
		Addr <=  "0010111000010";
		Trees_din <= x"bcff8904";
		wait for Clk_period;
		Addr <=  "0010111000011";
		Trees_din <= x"00a018d9";
		wait for Clk_period;
		Addr <=  "0010111000100";
		Trees_din <= x"ff9d18d9";
		wait for Clk_period;
		Addr <=  "0010111000101";
		Trees_din <= x"ff8e18d9";
		wait for Clk_period;
		Addr <=  "0010111000110";
		Trees_din <= x"1effc208";
		wait for Clk_period;
		Addr <=  "0010111000111";
		Trees_din <= x"39ff4b04";
		wait for Clk_period;
		Addr <=  "0010111001000";
		Trees_din <= x"ff8f18d9";
		wait for Clk_period;
		Addr <=  "0010111001001";
		Trees_din <= x"006f18d9";
		wait for Clk_period;
		Addr <=  "0010111001010";
		Trees_din <= x"08005604";
		wait for Clk_period;
		Addr <=  "0010111001011";
		Trees_din <= x"ff6918d9";
		wait for Clk_period;
		Addr <=  "0010111001100";
		Trees_din <= x"002f18d9";
		wait for Clk_period;
		Addr <=  "0010111001101";
		Trees_din <= x"03000f10";
		wait for Clk_period;
		Addr <=  "0010111001110";
		Trees_din <= x"27006b08";
		wait for Clk_period;
		Addr <=  "0010111001111";
		Trees_din <= x"b8fe9d04";
		wait for Clk_period;
		Addr <=  "0010111010000";
		Trees_din <= x"000418d9";
		wait for Clk_period;
		Addr <=  "0010111010001";
		Trees_din <= x"ff5e18d9";
		wait for Clk_period;
		Addr <=  "0010111010010";
		Trees_din <= x"97ff1104";
		wait for Clk_period;
		Addr <=  "0010111010011";
		Trees_din <= x"004c18d9";
		wait for Clk_period;
		Addr <=  "0010111010100";
		Trees_din <= x"000318d9";
		wait for Clk_period;
		Addr <=  "0010111010101";
		Trees_din <= x"e4fe9204";
		wait for Clk_period;
		Addr <=  "0010111010110";
		Trees_din <= x"ff9818d9";
		wait for Clk_period;
		Addr <=  "0010111010111";
		Trees_din <= x"3bff3604";
		wait for Clk_period;
		Addr <=  "0010111011000";
		Trees_din <= x"ffcb18d9";
		wait for Clk_period;
		Addr <=  "0010111011001";
		Trees_din <= x"00a118d9";
		wait for Clk_period;
		Addr <=  "0010111011010";
		Trees_din <= x"bcfee81c";
		wait for Clk_period;
		Addr <=  "0010111011011";
		Trees_din <= x"75ffdf0c";
		wait for Clk_period;
		Addr <=  "0010111011100";
		Trees_din <= x"77ffa108";
		wait for Clk_period;
		Addr <=  "0010111011101";
		Trees_din <= x"fb002f04";
		wait for Clk_period;
		Addr <=  "0010111011110";
		Trees_din <= x"008618d9";
		wait for Clk_period;
		Addr <=  "0010111011111";
		Trees_din <= x"ffaf18d9";
		wait for Clk_period;
		Addr <=  "0010111100000";
		Trees_din <= x"ff7c18d9";
		wait for Clk_period;
		Addr <=  "0010111100001";
		Trees_din <= x"d3ff5808";
		wait for Clk_period;
		Addr <=  "0010111100010";
		Trees_din <= x"74ffa004";
		wait for Clk_period;
		Addr <=  "0010111100011";
		Trees_din <= x"003d18d9";
		wait for Clk_period;
		Addr <=  "0010111100100";
		Trees_din <= x"ffc418d9";
		wait for Clk_period;
		Addr <=  "0010111100101";
		Trees_din <= x"3aff2604";
		wait for Clk_period;
		Addr <=  "0010111100110";
		Trees_din <= x"ffdc18d9";
		wait for Clk_period;
		Addr <=  "0010111100111";
		Trees_din <= x"00a418d9";
		wait for Clk_period;
		Addr <=  "0010111101000";
		Trees_din <= x"5c004110";
		wait for Clk_period;
		Addr <=  "0010111101001";
		Trees_din <= x"cafd9a08";
		wait for Clk_period;
		Addr <=  "0010111101010";
		Trees_din <= x"32fefa04";
		wait for Clk_period;
		Addr <=  "0010111101011";
		Trees_din <= x"ffc918d9";
		wait for Clk_period;
		Addr <=  "0010111101100";
		Trees_din <= x"00c018d9";
		wait for Clk_period;
		Addr <=  "0010111101101";
		Trees_din <= x"17007a04";
		wait for Clk_period;
		Addr <=  "0010111101110";
		Trees_din <= x"ffae18d9";
		wait for Clk_period;
		Addr <=  "0010111101111";
		Trees_din <= x"005718d9";
		wait for Clk_period;
		Addr <=  "0010111110000";
		Trees_din <= x"6f000908";
		wait for Clk_period;
		Addr <=  "0010111110001";
		Trees_din <= x"60ff7a04";
		wait for Clk_period;
		Addr <=  "0010111110010";
		Trees_din <= x"ffab18d9";
		wait for Clk_period;
		Addr <=  "0010111110011";
		Trees_din <= x"003318d9";
		wait for Clk_period;
		Addr <=  "0010111110100";
		Trees_din <= x"49ffef04";
		wait for Clk_period;
		Addr <=  "0010111110101";
		Trees_din <= x"002418d9";
		wait for Clk_period;
		Addr <=  "0010111110110";
		Trees_din <= x"00eb18d9";
		wait for Clk_period;
		Addr <=  "0010111110111";
		Trees_din <= x"28ff2e40";
		wait for Clk_period;
		Addr <=  "0010111111000";
		Trees_din <= x"f1ff9e20";
		wait for Clk_period;
		Addr <=  "0010111111001";
		Trees_din <= x"74000110";
		wait for Clk_period;
		Addr <=  "0010111111010";
		Trees_din <= x"8cff8d08";
		wait for Clk_period;
		Addr <=  "0010111111011";
		Trees_din <= x"8affa504";
		wait for Clk_period;
		Addr <=  "0010111111100";
		Trees_din <= x"005918d9";
		wait for Clk_period;
		Addr <=  "0010111111101";
		Trees_din <= x"ffb818d9";
		wait for Clk_period;
		Addr <=  "0010111111110";
		Trees_din <= x"8afef104";
		wait for Clk_period;
		Addr <=  "0010111111111";
		Trees_din <= x"ffe518d9";
		wait for Clk_period;
		Addr <=  "0011000000000";
		Trees_din <= x"008d18d9";
		wait for Clk_period;
		Addr <=  "0011000000001";
		Trees_din <= x"1eff8a08";
		wait for Clk_period;
		Addr <=  "0011000000010";
		Trees_din <= x"46ff4c04";
		wait for Clk_period;
		Addr <=  "0011000000011";
		Trees_din <= x"006118d9";
		wait for Clk_period;
		Addr <=  "0011000000100";
		Trees_din <= x"ff8518d9";
		wait for Clk_period;
		Addr <=  "0011000000101";
		Trees_din <= x"33fef204";
		wait for Clk_period;
		Addr <=  "0011000000110";
		Trees_din <= x"005718d9";
		wait for Clk_period;
		Addr <=  "0011000000111";
		Trees_din <= x"ff8d18d9";
		wait for Clk_period;
		Addr <=  "0011000001000";
		Trees_din <= x"ee003710";
		wait for Clk_period;
		Addr <=  "0011000001001";
		Trees_din <= x"30001a08";
		wait for Clk_period;
		Addr <=  "0011000001010";
		Trees_din <= x"c5ff8404";
		wait for Clk_period;
		Addr <=  "0011000001011";
		Trees_din <= x"004f18d9";
		wait for Clk_period;
		Addr <=  "0011000001100";
		Trees_din <= x"ffa318d9";
		wait for Clk_period;
		Addr <=  "0011000001101";
		Trees_din <= x"91ff2804";
		wait for Clk_period;
		Addr <=  "0011000001110";
		Trees_din <= x"004718d9";
		wait for Clk_period;
		Addr <=  "0011000001111";
		Trees_din <= x"ff8918d9";
		wait for Clk_period;
		Addr <=  "0011000010000";
		Trees_din <= x"26006008";
		wait for Clk_period;
		Addr <=  "0011000010001";
		Trees_din <= x"f5008104";
		wait for Clk_period;
		Addr <=  "0011000010010";
		Trees_din <= x"ff6518d9";
		wait for Clk_period;
		Addr <=  "0011000010011";
		Trees_din <= x"006918d9";
		wait for Clk_period;
		Addr <=  "0011000010100";
		Trees_din <= x"c3fff504";
		wait for Clk_period;
		Addr <=  "0011000010101";
		Trees_din <= x"ffbb18d9";
		wait for Clk_period;
		Addr <=  "0011000010110";
		Trees_din <= x"005718d9";
		wait for Clk_period;
		Addr <=  "0011000010111";
		Trees_din <= x"61ff6820";
		wait for Clk_period;
		Addr <=  "0011000011000";
		Trees_din <= x"ab004310";
		wait for Clk_period;
		Addr <=  "0011000011001";
		Trees_din <= x"05003208";
		wait for Clk_period;
		Addr <=  "0011000011010";
		Trees_din <= x"61fe7304";
		wait for Clk_period;
		Addr <=  "0011000011011";
		Trees_din <= x"006618d9";
		wait for Clk_period;
		Addr <=  "0011000011100";
		Trees_din <= x"ff6f18d9";
		wait for Clk_period;
		Addr <=  "0011000011101";
		Trees_din <= x"afff1f04";
		wait for Clk_period;
		Addr <=  "0011000011110";
		Trees_din <= x"ff9d18d9";
		wait for Clk_period;
		Addr <=  "0011000011111";
		Trees_din <= x"005518d9";
		wait for Clk_period;
		Addr <=  "0011000100000";
		Trees_din <= x"a0feaa08";
		wait for Clk_period;
		Addr <=  "0011000100001";
		Trees_din <= x"3eff9a04";
		wait for Clk_period;
		Addr <=  "0011000100010";
		Trees_din <= x"ffc018d9";
		wait for Clk_period;
		Addr <=  "0011000100011";
		Trees_din <= x"007618d9";
		wait for Clk_period;
		Addr <=  "0011000100100";
		Trees_din <= x"8e00e604";
		wait for Clk_period;
		Addr <=  "0011000100101";
		Trees_din <= x"ff7618d9";
		wait for Clk_period;
		Addr <=  "0011000100110";
		Trees_din <= x"007518d9";
		wait for Clk_period;
		Addr <=  "0011000100111";
		Trees_din <= x"89004710";
		wait for Clk_period;
		Addr <=  "0011000101000";
		Trees_din <= x"5a003e08";
		wait for Clk_period;
		Addr <=  "0011000101001";
		Trees_din <= x"27ffc504";
		wait for Clk_period;
		Addr <=  "0011000101010";
		Trees_din <= x"ffa418d9";
		wait for Clk_period;
		Addr <=  "0011000101011";
		Trees_din <= x"003918d9";
		wait for Clk_period;
		Addr <=  "0011000101100";
		Trees_din <= x"a7ff3804";
		wait for Clk_period;
		Addr <=  "0011000101101";
		Trees_din <= x"fff118d9";
		wait for Clk_period;
		Addr <=  "0011000101110";
		Trees_din <= x"006318d9";
		wait for Clk_period;
		Addr <=  "0011000101111";
		Trees_din <= x"58fea608";
		wait for Clk_period;
		Addr <=  "0011000110000";
		Trees_din <= x"bbffa004";
		wait for Clk_period;
		Addr <=  "0011000110001";
		Trees_din <= x"ffd118d9";
		wait for Clk_period;
		Addr <=  "0011000110010";
		Trees_din <= x"00c918d9";
		wait for Clk_period;
		Addr <=  "0011000110011";
		Trees_din <= x"f4ff5a04";
		wait for Clk_period;
		Addr <=  "0011000110100";
		Trees_din <= x"ff5818d9";
		wait for Clk_period;
		Addr <=  "0011000110101";
		Trees_din <= x"007018d9";
		wait for Clk_period;
		Addr <=  "0011000110110";
		Trees_din <= x"36fee954";
		wait for Clk_period;
		Addr <=  "0011000110111";
		Trees_din <= x"b8ff1630";
		wait for Clk_period;
		Addr <=  "0011000111000";
		Trees_din <= x"85ff9a14";
		wait for Clk_period;
		Addr <=  "0011000111001";
		Trees_din <= x"19ff3408";
		wait for Clk_period;
		Addr <=  "0011000111010";
		Trees_din <= x"33fece04";
		wait for Clk_period;
		Addr <=  "0011000111011";
		Trees_din <= x"007c1a4d";
		wait for Clk_period;
		Addr <=  "0011000111100";
		Trees_din <= x"ff961a4d";
		wait for Clk_period;
		Addr <=  "0011000111101";
		Trees_din <= x"0fffc908";
		wait for Clk_period;
		Addr <=  "0011000111110";
		Trees_din <= x"0fff3604";
		wait for Clk_period;
		Addr <=  "0011000111111";
		Trees_din <= x"001d1a4d";
		wait for Clk_period;
		Addr <=  "0011001000000";
		Trees_din <= x"00e21a4d";
		wait for Clk_period;
		Addr <=  "0011001000001";
		Trees_din <= x"fff01a4d";
		wait for Clk_period;
		Addr <=  "0011001000010";
		Trees_din <= x"4bfe7a0c";
		wait for Clk_period;
		Addr <=  "0011001000011";
		Trees_din <= x"61ffb308";
		wait for Clk_period;
		Addr <=  "0011001000100";
		Trees_din <= x"0dff8204";
		wait for Clk_period;
		Addr <=  "0011001000101";
		Trees_din <= x"00b31a4d";
		wait for Clk_period;
		Addr <=  "0011001000110";
		Trees_din <= x"000b1a4d";
		wait for Clk_period;
		Addr <=  "0011001000111";
		Trees_din <= x"ffa71a4d";
		wait for Clk_period;
		Addr <=  "0011001001000";
		Trees_din <= x"a0ff3208";
		wait for Clk_period;
		Addr <=  "0011001001001";
		Trees_din <= x"19ff0604";
		wait for Clk_period;
		Addr <=  "0011001001010";
		Trees_din <= x"fff61a4d";
		wait for Clk_period;
		Addr <=  "0011001001011";
		Trees_din <= x"ff691a4d";
		wait for Clk_period;
		Addr <=  "0011001001100";
		Trees_din <= x"f4ff0004";
		wait for Clk_period;
		Addr <=  "0011001001101";
		Trees_din <= x"00701a4d";
		wait for Clk_period;
		Addr <=  "0011001001110";
		Trees_din <= x"ffb01a4d";
		wait for Clk_period;
		Addr <=  "0011001001111";
		Trees_din <= x"e8fe6604";
		wait for Clk_period;
		Addr <=  "0011001010000";
		Trees_din <= x"00b11a4d";
		wait for Clk_period;
		Addr <=  "0011001010001";
		Trees_din <= x"86fe8810";
		wait for Clk_period;
		Addr <=  "0011001010010";
		Trees_din <= x"54005308";
		wait for Clk_period;
		Addr <=  "0011001010011";
		Trees_din <= x"d1ff0104";
		wait for Clk_period;
		Addr <=  "0011001010100";
		Trees_din <= x"00461a4d";
		wait for Clk_period;
		Addr <=  "0011001010101";
		Trees_din <= x"ff771a4d";
		wait for Clk_period;
		Addr <=  "0011001010110";
		Trees_din <= x"04005104";
		wait for Clk_period;
		Addr <=  "0011001010111";
		Trees_din <= x"ffba1a4d";
		wait for Clk_period;
		Addr <=  "0011001011000";
		Trees_din <= x"00951a4d";
		wait for Clk_period;
		Addr <=  "0011001011001";
		Trees_din <= x"0ffff008";
		wait for Clk_period;
		Addr <=  "0011001011010";
		Trees_din <= x"0effa904";
		wait for Clk_period;
		Addr <=  "0011001011011";
		Trees_din <= x"ff8c1a4d";
		wait for Clk_period;
		Addr <=  "0011001011100";
		Trees_din <= x"00731a4d";
		wait for Clk_period;
		Addr <=  "0011001011101";
		Trees_din <= x"faff9f04";
		wait for Clk_period;
		Addr <=  "0011001011110";
		Trees_din <= x"ffc71a4d";
		wait for Clk_period;
		Addr <=  "0011001011111";
		Trees_din <= x"00a11a4d";
		wait for Clk_period;
		Addr <=  "0011001100000";
		Trees_din <= x"5dffe13c";
		wait for Clk_period;
		Addr <=  "0011001100001";
		Trees_din <= x"a5feb41c";
		wait for Clk_period;
		Addr <=  "0011001100010";
		Trees_din <= x"34004310";
		wait for Clk_period;
		Addr <=  "0011001100011";
		Trees_din <= x"2eff3508";
		wait for Clk_period;
		Addr <=  "0011001100100";
		Trees_din <= x"99fef104";
		wait for Clk_period;
		Addr <=  "0011001100101";
		Trees_din <= x"009e1a4d";
		wait for Clk_period;
		Addr <=  "0011001100110";
		Trees_din <= x"ff9d1a4d";
		wait for Clk_period;
		Addr <=  "0011001100111";
		Trees_din <= x"cc006404";
		wait for Clk_period;
		Addr <=  "0011001101000";
		Trees_din <= x"ff901a4d";
		wait for Clk_period;
		Addr <=  "0011001101001";
		Trees_din <= x"00351a4d";
		wait for Clk_period;
		Addr <=  "0011001101010";
		Trees_din <= x"8effa704";
		wait for Clk_period;
		Addr <=  "0011001101011";
		Trees_din <= x"ff931a4d";
		wait for Clk_period;
		Addr <=  "0011001101100";
		Trees_din <= x"8e004f04";
		wait for Clk_period;
		Addr <=  "0011001101101";
		Trees_din <= x"00d31a4d";
		wait for Clk_period;
		Addr <=  "0011001101110";
		Trees_din <= x"ffc71a4d";
		wait for Clk_period;
		Addr <=  "0011001101111";
		Trees_din <= x"cffffd10";
		wait for Clk_period;
		Addr <=  "0011001110000";
		Trees_din <= x"00ff5208";
		wait for Clk_period;
		Addr <=  "0011001110001";
		Trees_din <= x"d7ffe504";
		wait for Clk_period;
		Addr <=  "0011001110010";
		Trees_din <= x"ff751a4d";
		wait for Clk_period;
		Addr <=  "0011001110011";
		Trees_din <= x"00401a4d";
		wait for Clk_period;
		Addr <=  "0011001110100";
		Trees_din <= x"6ffff904";
		wait for Clk_period;
		Addr <=  "0011001110101";
		Trees_din <= x"ffc61a4d";
		wait for Clk_period;
		Addr <=  "0011001110110";
		Trees_din <= x"00631a4d";
		wait for Clk_period;
		Addr <=  "0011001110111";
		Trees_din <= x"3eff9508";
		wait for Clk_period;
		Addr <=  "0011001111000";
		Trees_din <= x"30000c04";
		wait for Clk_period;
		Addr <=  "0011001111001";
		Trees_din <= x"00351a4d";
		wait for Clk_period;
		Addr <=  "0011001111010";
		Trees_din <= x"ffef1a4d";
		wait for Clk_period;
		Addr <=  "0011001111011";
		Trees_din <= x"1cff5004";
		wait for Clk_period;
		Addr <=  "0011001111100";
		Trees_din <= x"00321a4d";
		wait for Clk_period;
		Addr <=  "0011001111101";
		Trees_din <= x"008a1a4d";
		wait for Clk_period;
		Addr <=  "0011001111110";
		Trees_din <= x"3b004520";
		wait for Clk_period;
		Addr <=  "0011001111111";
		Trees_din <= x"ceffe710";
		wait for Clk_period;
		Addr <=  "0011010000000";
		Trees_din <= x"83ffc608";
		wait for Clk_period;
		Addr <=  "0011010000001";
		Trees_din <= x"c3ffdc04";
		wait for Clk_period;
		Addr <=  "0011010000010";
		Trees_din <= x"ffa51a4d";
		wait for Clk_period;
		Addr <=  "0011010000011";
		Trees_din <= x"fff21a4d";
		wait for Clk_period;
		Addr <=  "0011010000100";
		Trees_din <= x"46feba04";
		wait for Clk_period;
		Addr <=  "0011010000101";
		Trees_din <= x"00d91a4d";
		wait for Clk_period;
		Addr <=  "0011010000110";
		Trees_din <= x"000b1a4d";
		wait for Clk_period;
		Addr <=  "0011010000111";
		Trees_din <= x"c2ff7308";
		wait for Clk_period;
		Addr <=  "0011010001000";
		Trees_din <= x"40fff804";
		wait for Clk_period;
		Addr <=  "0011010001001";
		Trees_din <= x"ff8a1a4d";
		wait for Clk_period;
		Addr <=  "0011010001010";
		Trees_din <= x"001a1a4d";
		wait for Clk_period;
		Addr <=  "0011010001011";
		Trees_din <= x"f3ff6e04";
		wait for Clk_period;
		Addr <=  "0011010001100";
		Trees_din <= x"005f1a4d";
		wait for Clk_period;
		Addr <=  "0011010001101";
		Trees_din <= x"ff991a4d";
		wait for Clk_period;
		Addr <=  "0011010001110";
		Trees_din <= x"0cfe4d04";
		wait for Clk_period;
		Addr <=  "0011010001111";
		Trees_din <= x"ffe41a4d";
		wait for Clk_period;
		Addr <=  "0011010010000";
		Trees_din <= x"e6ff5104";
		wait for Clk_period;
		Addr <=  "0011010010001";
		Trees_din <= x"00351a4d";
		wait for Clk_period;
		Addr <=  "0011010010010";
		Trees_din <= x"00e91a4d";
		wait for Clk_period;
		Addr <=  "0011010010011";
		Trees_din <= x"09001e78";
		wait for Clk_period;
		Addr <=  "0011010010100";
		Trees_din <= x"43ffa740";
		wait for Clk_period;
		Addr <=  "0011010010101";
		Trees_din <= x"87ff7b20";
		wait for Clk_period;
		Addr <=  "0011010010110";
		Trees_din <= x"04ffc210";
		wait for Clk_period;
		Addr <=  "0011010010111";
		Trees_din <= x"98ff6b08";
		wait for Clk_period;
		Addr <=  "0011010011000";
		Trees_din <= x"3bffe604";
		wait for Clk_period;
		Addr <=  "0011010011001";
		Trees_din <= x"ff641bb9";
		wait for Clk_period;
		Addr <=  "0011010011010";
		Trees_din <= x"002f1bb9";
		wait for Clk_period;
		Addr <=  "0011010011011";
		Trees_din <= x"1bff9504";
		wait for Clk_period;
		Addr <=  "0011010011100";
		Trees_din <= x"ffd61bb9";
		wait for Clk_period;
		Addr <=  "0011010011101";
		Trees_din <= x"00ad1bb9";
		wait for Clk_period;
		Addr <=  "0011010011110";
		Trees_din <= x"11fff008";
		wait for Clk_period;
		Addr <=  "0011010011111";
		Trees_din <= x"ec001904";
		wait for Clk_period;
		Addr <=  "0011010100000";
		Trees_din <= x"00171bb9";
		wait for Clk_period;
		Addr <=  "0011010100001";
		Trees_din <= x"004c1bb9";
		wait for Clk_period;
		Addr <=  "0011010100010";
		Trees_din <= x"34005304";
		wait for Clk_period;
		Addr <=  "0011010100011";
		Trees_din <= x"ff9a1bb9";
		wait for Clk_period;
		Addr <=  "0011010100100";
		Trees_din <= x"00711bb9";
		wait for Clk_period;
		Addr <=  "0011010100101";
		Trees_din <= x"1effbd10";
		wait for Clk_period;
		Addr <=  "0011010100110";
		Trees_din <= x"a0fe0408";
		wait for Clk_period;
		Addr <=  "0011010100111";
		Trees_din <= x"8aff0504";
		wait for Clk_period;
		Addr <=  "0011010101000";
		Trees_din <= x"00501bb9";
		wait for Clk_period;
		Addr <=  "0011010101001";
		Trees_din <= x"ff561bb9";
		wait for Clk_period;
		Addr <=  "0011010101010";
		Trees_din <= x"d9ff9004";
		wait for Clk_period;
		Addr <=  "0011010101011";
		Trees_din <= x"004d1bb9";
		wait for Clk_period;
		Addr <=  "0011010101100";
		Trees_din <= x"fffa1bb9";
		wait for Clk_period;
		Addr <=  "0011010101101";
		Trees_din <= x"f1ff8b08";
		wait for Clk_period;
		Addr <=  "0011010101110";
		Trees_din <= x"38ff8104";
		wait for Clk_period;
		Addr <=  "0011010101111";
		Trees_din <= x"003c1bb9";
		wait for Clk_period;
		Addr <=  "0011010110000";
		Trees_din <= x"ff921bb9";
		wait for Clk_period;
		Addr <=  "0011010110001";
		Trees_din <= x"90fed204";
		wait for Clk_period;
		Addr <=  "0011010110010";
		Trees_din <= x"002e1bb9";
		wait for Clk_period;
		Addr <=  "0011010110011";
		Trees_din <= x"ff851bb9";
		wait for Clk_period;
		Addr <=  "0011010110100";
		Trees_din <= x"16fe3918";
		wait for Clk_period;
		Addr <=  "0011010110101";
		Trees_din <= x"00ff460c";
		wait for Clk_period;
		Addr <=  "0011010110110";
		Trees_din <= x"e4fe1904";
		wait for Clk_period;
		Addr <=  "0011010110111";
		Trees_din <= x"ffc11bb9";
		wait for Clk_period;
		Addr <=  "0011010111000";
		Trees_din <= x"85ffe404";
		wait for Clk_period;
		Addr <=  "0011010111001";
		Trees_din <= x"00f21bb9";
		wait for Clk_period;
		Addr <=  "0011010111010";
		Trees_din <= x"fff91bb9";
		wait for Clk_period;
		Addr <=  "0011010111011";
		Trees_din <= x"53ffec08";
		wait for Clk_period;
		Addr <=  "0011010111100";
		Trees_din <= x"69ff1104";
		wait for Clk_period;
		Addr <=  "0011010111101";
		Trees_din <= x"ffe81bb9";
		wait for Clk_period;
		Addr <=  "0011010111110";
		Trees_din <= x"ff7f1bb9";
		wait for Clk_period;
		Addr <=  "0011010111111";
		Trees_din <= x"00601bb9";
		wait for Clk_period;
		Addr <=  "0011011000000";
		Trees_din <= x"31005210";
		wait for Clk_period;
		Addr <=  "0011011000001";
		Trees_din <= x"33ff2b08";
		wait for Clk_period;
		Addr <=  "0011011000010";
		Trees_din <= x"67ffa804";
		wait for Clk_period;
		Addr <=  "0011011000011";
		Trees_din <= x"ffc81bb9";
		wait for Clk_period;
		Addr <=  "0011011000100";
		Trees_din <= x"004c1bb9";
		wait for Clk_period;
		Addr <=  "0011011000101";
		Trees_din <= x"0a00e004";
		wait for Clk_period;
		Addr <=  "0011011000110";
		Trees_din <= x"ff821bb9";
		wait for Clk_period;
		Addr <=  "0011011000111";
		Trees_din <= x"003e1bb9";
		wait for Clk_period;
		Addr <=  "0011011001000";
		Trees_din <= x"74ffd308";
		wait for Clk_period;
		Addr <=  "0011011001001";
		Trees_din <= x"c1fe9304";
		wait for Clk_period;
		Addr <=  "0011011001010";
		Trees_din <= x"00561bb9";
		wait for Clk_period;
		Addr <=  "0011011001011";
		Trees_din <= x"ff751bb9";
		wait for Clk_period;
		Addr <=  "0011011001100";
		Trees_din <= x"3cff2204";
		wait for Clk_period;
		Addr <=  "0011011001101";
		Trees_din <= x"008f1bb9";
		wait for Clk_period;
		Addr <=  "0011011001110";
		Trees_din <= x"ffa11bb9";
		wait for Clk_period;
		Addr <=  "0011011001111";
		Trees_din <= x"39ff1f0c";
		wait for Clk_period;
		Addr <=  "0011011010000";
		Trees_din <= x"60ffec08";
		wait for Clk_period;
		Addr <=  "0011011010001";
		Trees_din <= x"b2ff5b04";
		wait for Clk_period;
		Addr <=  "0011011010010";
		Trees_din <= x"ffdd1bb9";
		wait for Clk_period;
		Addr <=  "0011011010011";
		Trees_din <= x"ff621bb9";
		wait for Clk_period;
		Addr <=  "0011011010100";
		Trees_din <= x"007e1bb9";
		wait for Clk_period;
		Addr <=  "0011011010101";
		Trees_din <= x"85ff0814";
		wait for Clk_period;
		Addr <=  "0011011010110";
		Trees_din <= x"15ffc70c";
		wait for Clk_period;
		Addr <=  "0011011010111";
		Trees_din <= x"21ff2c04";
		wait for Clk_period;
		Addr <=  "0011011011000";
		Trees_din <= x"ffc41bb9";
		wait for Clk_period;
		Addr <=  "0011011011001";
		Trees_din <= x"58fe2904";
		wait for Clk_period;
		Addr <=  "0011011011010";
		Trees_din <= x"ffe61bb9";
		wait for Clk_period;
		Addr <=  "0011011011011";
		Trees_din <= x"00c01bb9";
		wait for Clk_period;
		Addr <=  "0011011011100";
		Trees_din <= x"91ff8004";
		wait for Clk_period;
		Addr <=  "0011011011101";
		Trees_din <= x"ff891bb9";
		wait for Clk_period;
		Addr <=  "0011011011110";
		Trees_din <= x"00821bb9";
		wait for Clk_period;
		Addr <=  "0011011011111";
		Trees_din <= x"97ff1510";
		wait for Clk_period;
		Addr <=  "0011011100000";
		Trees_din <= x"f8006808";
		wait for Clk_period;
		Addr <=  "0011011100001";
		Trees_din <= x"80ff5304";
		wait for Clk_period;
		Addr <=  "0011011100010";
		Trees_din <= x"00771bb9";
		wait for Clk_period;
		Addr <=  "0011011100011";
		Trees_din <= x"ffed1bb9";
		wait for Clk_period;
		Addr <=  "0011011100100";
		Trees_din <= x"7bff6904";
		wait for Clk_period;
		Addr <=  "0011011100101";
		Trees_din <= x"ff721bb9";
		wait for Clk_period;
		Addr <=  "0011011100110";
		Trees_din <= x"002e1bb9";
		wait for Clk_period;
		Addr <=  "0011011100111";
		Trees_din <= x"bdffcf08";
		wait for Clk_period;
		Addr <=  "0011011101000";
		Trees_din <= x"2fffa904";
		wait for Clk_period;
		Addr <=  "0011011101001";
		Trees_din <= x"ffdb1bb9";
		wait for Clk_period;
		Addr <=  "0011011101010";
		Trees_din <= x"00611bb9";
		wait for Clk_period;
		Addr <=  "0011011101011";
		Trees_din <= x"4eff6b04";
		wait for Clk_period;
		Addr <=  "0011011101100";
		Trees_din <= x"00a91bb9";
		wait for Clk_period;
		Addr <=  "0011011101101";
		Trees_din <= x"00381bb9";
		wait for Clk_period;
		Addr <=  "0011011101110";
		Trees_din <= x"3d00277c";
		wait for Clk_period;
		Addr <=  "0011011101111";
		Trees_din <= x"25007840";
		wait for Clk_period;
		Addr <=  "0011011110000";
		Trees_din <= x"36ffcb20";
		wait for Clk_period;
		Addr <=  "0011011110001";
		Trees_din <= x"8aff9b10";
		wait for Clk_period;
		Addr <=  "0011011110010";
		Trees_din <= x"0efe3508";
		wait for Clk_period;
		Addr <=  "0011011110011";
		Trees_din <= x"fbffab04";
		wait for Clk_period;
		Addr <=  "0011011110100";
		Trees_din <= x"001a1d5d";
		wait for Clk_period;
		Addr <=  "0011011110101";
		Trees_din <= x"009b1d5d";
		wait for Clk_period;
		Addr <=  "0011011110110";
		Trees_din <= x"95fed804";
		wait for Clk_period;
		Addr <=  "0011011110111";
		Trees_din <= x"00441d5d";
		wait for Clk_period;
		Addr <=  "0011011111000";
		Trees_din <= x"fff61d5d";
		wait for Clk_period;
		Addr <=  "0011011111001";
		Trees_din <= x"ebfea908";
		wait for Clk_period;
		Addr <=  "0011011111010";
		Trees_din <= x"4dfe6804";
		wait for Clk_period;
		Addr <=  "0011011111011";
		Trees_din <= x"005f1d5d";
		wait for Clk_period;
		Addr <=  "0011011111100";
		Trees_din <= x"fff21d5d";
		wait for Clk_period;
		Addr <=  "0011011111101";
		Trees_din <= x"41ff5904";
		wait for Clk_period;
		Addr <=  "0011011111110";
		Trees_din <= x"ffe41d5d";
		wait for Clk_period;
		Addr <=  "0011011111111";
		Trees_din <= x"ff891d5d";
		wait for Clk_period;
		Addr <=  "0011100000000";
		Trees_din <= x"73fff410";
		wait for Clk_period;
		Addr <=  "0011100000001";
		Trees_din <= x"74ffe908";
		wait for Clk_period;
		Addr <=  "0011100000010";
		Trees_din <= x"bfff9404";
		wait for Clk_period;
		Addr <=  "0011100000011";
		Trees_din <= x"008d1d5d";
		wait for Clk_period;
		Addr <=  "0011100000100";
		Trees_din <= x"ffba1d5d";
		wait for Clk_period;
		Addr <=  "0011100000101";
		Trees_din <= x"cc003904";
		wait for Clk_period;
		Addr <=  "0011100000110";
		Trees_din <= x"ffa01d5d";
		wait for Clk_period;
		Addr <=  "0011100000111";
		Trees_din <= x"003f1d5d";
		wait for Clk_period;
		Addr <=  "0011100001000";
		Trees_din <= x"f4fe8108";
		wait for Clk_period;
		Addr <=  "0011100001001";
		Trees_din <= x"21ff8e04";
		wait for Clk_period;
		Addr <=  "0011100001010";
		Trees_din <= x"00681d5d";
		wait for Clk_period;
		Addr <=  "0011100001011";
		Trees_din <= x"ff9b1d5d";
		wait for Clk_period;
		Addr <=  "0011100001100";
		Trees_din <= x"29ffda04";
		wait for Clk_period;
		Addr <=  "0011100001101";
		Trees_din <= x"00af1d5d";
		wait for Clk_period;
		Addr <=  "0011100001110";
		Trees_din <= x"fff01d5d";
		wait for Clk_period;
		Addr <=  "0011100001111";
		Trees_din <= x"00ff961c";
		wait for Clk_period;
		Addr <=  "0011100010000";
		Trees_din <= x"bcff190c";
		wait for Clk_period;
		Addr <=  "0011100010001";
		Trees_din <= x"21006008";
		wait for Clk_period;
		Addr <=  "0011100010010";
		Trees_din <= x"e6003204";
		wait for Clk_period;
		Addr <=  "0011100010011";
		Trees_din <= x"007e1d5d";
		wait for Clk_period;
		Addr <=  "0011100010100";
		Trees_din <= x"ffbe1d5d";
		wait for Clk_period;
		Addr <=  "0011100010101";
		Trees_din <= x"ff791d5d";
		wait for Clk_period;
		Addr <=  "0011100010110";
		Trees_din <= x"e5fee408";
		wait for Clk_period;
		Addr <=  "0011100010111";
		Trees_din <= x"46feb304";
		wait for Clk_period;
		Addr <=  "0011100011000";
		Trees_din <= x"ffb31d5d";
		wait for Clk_period;
		Addr <=  "0011100011001";
		Trees_din <= x"00681d5d";
		wait for Clk_period;
		Addr <=  "0011100011010";
		Trees_din <= x"88fff404";
		wait for Clk_period;
		Addr <=  "0011100011011";
		Trees_din <= x"002e1d5d";
		wait for Clk_period;
		Addr <=  "0011100011100";
		Trees_din <= x"ff811d5d";
		wait for Clk_period;
		Addr <=  "0011100011101";
		Trees_din <= x"33ff0a10";
		wait for Clk_period;
		Addr <=  "0011100011110";
		Trees_din <= x"24ff2a08";
		wait for Clk_period;
		Addr <=  "0011100011111";
		Trees_din <= x"22ff8c04";
		wait for Clk_period;
		Addr <=  "0011100100000";
		Trees_din <= x"ffec1d5d";
		wait for Clk_period;
		Addr <=  "0011100100001";
		Trees_din <= x"ff7e1d5d";
		wait for Clk_period;
		Addr <=  "0011100100010";
		Trees_din <= x"00001d04";
		wait for Clk_period;
		Addr <=  "0011100100011";
		Trees_din <= x"008f1d5d";
		wait for Clk_period;
		Addr <=  "0011100100100";
		Trees_din <= x"ff961d5d";
		wait for Clk_period;
		Addr <=  "0011100100101";
		Trees_din <= x"8e003b08";
		wait for Clk_period;
		Addr <=  "0011100100110";
		Trees_din <= x"d5005704";
		wait for Clk_period;
		Addr <=  "0011100100111";
		Trees_din <= x"ff651d5d";
		wait for Clk_period;
		Addr <=  "0011100101000";
		Trees_din <= x"00351d5d";
		wait for Clk_period;
		Addr <=  "0011100101001";
		Trees_din <= x"f8001004";
		wait for Clk_period;
		Addr <=  "0011100101010";
		Trees_din <= x"008e1d5d";
		wait for Clk_period;
		Addr <=  "0011100101011";
		Trees_din <= x"ffe41d5d";
		wait for Clk_period;
		Addr <=  "0011100101100";
		Trees_din <= x"e0fe7220";
		wait for Clk_period;
		Addr <=  "0011100101101";
		Trees_din <= x"9eff4b10";
		wait for Clk_period;
		Addr <=  "0011100101110";
		Trees_din <= x"9fff0108";
		wait for Clk_period;
		Addr <=  "0011100101111";
		Trees_din <= x"18ff8f04";
		wait for Clk_period;
		Addr <=  "0011100110000";
		Trees_din <= x"00831d5d";
		wait for Clk_period;
		Addr <=  "0011100110001";
		Trees_din <= x"00141d5d";
		wait for Clk_period;
		Addr <=  "0011100110010";
		Trees_din <= x"18fffb04";
		wait for Clk_period;
		Addr <=  "0011100110011";
		Trees_din <= x"ff761d5d";
		wait for Clk_period;
		Addr <=  "0011100110100";
		Trees_din <= x"00621d5d";
		wait for Clk_period;
		Addr <=  "0011100110101";
		Trees_din <= x"4eff980c";
		wait for Clk_period;
		Addr <=  "0011100110110";
		Trees_din <= x"06ff4004";
		wait for Clk_period;
		Addr <=  "0011100110111";
		Trees_din <= x"ffe11d5d";
		wait for Clk_period;
		Addr <=  "0011100111000";
		Trees_din <= x"71fe8804";
		wait for Clk_period;
		Addr <=  "0011100111001";
		Trees_din <= x"001d1d5d";
		wait for Clk_period;
		Addr <=  "0011100111010";
		Trees_din <= x"00e81d5d";
		wait for Clk_period;
		Addr <=  "0011100111011";
		Trees_din <= x"ffa21d5d";
		wait for Clk_period;
		Addr <=  "0011100111100";
		Trees_din <= x"7affa018";
		wait for Clk_period;
		Addr <=  "0011100111101";
		Trees_din <= x"71000210";
		wait for Clk_period;
		Addr <=  "0011100111110";
		Trees_din <= x"33ff0708";
		wait for Clk_period;
		Addr <=  "0011100111111";
		Trees_din <= x"99fefb04";
		wait for Clk_period;
		Addr <=  "0011101000000";
		Trees_din <= x"ffa51d5d";
		wait for Clk_period;
		Addr <=  "0011101000001";
		Trees_din <= x"002f1d5d";
		wait for Clk_period;
		Addr <=  "0011101000010";
		Trees_din <= x"a1fe9504";
		wait for Clk_period;
		Addr <=  "0011101000011";
		Trees_din <= x"fffc1d5d";
		wait for Clk_period;
		Addr <=  "0011101000100";
		Trees_din <= x"ff6e1d5d";
		wait for Clk_period;
		Addr <=  "0011101000101";
		Trees_din <= x"eeffe404";
		wait for Clk_period;
		Addr <=  "0011101000110";
		Trees_din <= x"ffd91d5d";
		wait for Clk_period;
		Addr <=  "0011101000111";
		Trees_din <= x"00d31d5d";
		wait for Clk_period;
		Addr <=  "0011101001000";
		Trees_din <= x"56ff7d10";
		wait for Clk_period;
		Addr <=  "0011101001001";
		Trees_din <= x"d8005f08";
		wait for Clk_period;
		Addr <=  "0011101001010";
		Trees_din <= x"fdfed104";
		wait for Clk_period;
		Addr <=  "0011101001011";
		Trees_din <= x"00531d5d";
		wait for Clk_period;
		Addr <=  "0011101001100";
		Trees_din <= x"ff8f1d5d";
		wait for Clk_period;
		Addr <=  "0011101001101";
		Trees_din <= x"88001304";
		wait for Clk_period;
		Addr <=  "0011101001110";
		Trees_din <= x"007d1d5d";
		wait for Clk_period;
		Addr <=  "0011101001111";
		Trees_din <= x"ffcf1d5d";
		wait for Clk_period;
		Addr <=  "0011101010000";
		Trees_din <= x"b9fed408";
		wait for Clk_period;
		Addr <=  "0011101010001";
		Trees_din <= x"95ff0c04";
		wait for Clk_period;
		Addr <=  "0011101010010";
		Trees_din <= x"00251d5d";
		wait for Clk_period;
		Addr <=  "0011101010011";
		Trees_din <= x"ff781d5d";
		wait for Clk_period;
		Addr <=  "0011101010100";
		Trees_din <= x"c7fef804";
		wait for Clk_period;
		Addr <=  "0011101010101";
		Trees_din <= x"00781d5d";
		wait for Clk_period;
		Addr <=  "0011101010110";
		Trees_din <= x"fff91d5d";
		wait for Clk_period;
		Addr <=  "0011101010111";
		Trees_din <= x"83ffc380";
		wait for Clk_period;
		Addr <=  "0011101011000";
		Trees_din <= x"7aff6640";
		wait for Clk_period;
		Addr <=  "0011101011001";
		Trees_din <= x"f4ff0820";
		wait for Clk_period;
		Addr <=  "0011101011010";
		Trees_din <= x"9ffefd10";
		wait for Clk_period;
		Addr <=  "0011101011011";
		Trees_din <= x"59fffd08";
		wait for Clk_period;
		Addr <=  "0011101011100";
		Trees_din <= x"30ffff04";
		wait for Clk_period;
		Addr <=  "0011101011101";
		Trees_din <= x"00a71f11";
		wait for Clk_period;
		Addr <=  "0011101011110";
		Trees_din <= x"fff61f11";
		wait for Clk_period;
		Addr <=  "0011101011111";
		Trees_din <= x"38fee004";
		wait for Clk_period;
		Addr <=  "0011101100000";
		Trees_din <= x"006f1f11";
		wait for Clk_period;
		Addr <=  "0011101100001";
		Trees_din <= x"ff7c1f11";
		wait for Clk_period;
		Addr <=  "0011101100010";
		Trees_din <= x"6d000308";
		wait for Clk_period;
		Addr <=  "0011101100011";
		Trees_din <= x"de007a04";
		wait for Clk_period;
		Addr <=  "0011101100100";
		Trees_din <= x"ff881f11";
		wait for Clk_period;
		Addr <=  "0011101100101";
		Trees_din <= x"002a1f11";
		wait for Clk_period;
		Addr <=  "0011101100110";
		Trees_din <= x"65ff7904";
		wait for Clk_period;
		Addr <=  "0011101100111";
		Trees_din <= x"00301f11";
		wait for Clk_period;
		Addr <=  "0011101101000";
		Trees_din <= x"ffb41f11";
		wait for Clk_period;
		Addr <=  "0011101101001";
		Trees_din <= x"bbff0f10";
		wait for Clk_period;
		Addr <=  "0011101101010";
		Trees_din <= x"39005e08";
		wait for Clk_period;
		Addr <=  "0011101101011";
		Trees_din <= x"42fed504";
		wait for Clk_period;
		Addr <=  "0011101101100";
		Trees_din <= x"001a1f11";
		wait for Clk_period;
		Addr <=  "0011101101101";
		Trees_din <= x"ff631f11";
		wait for Clk_period;
		Addr <=  "0011101101110";
		Trees_din <= x"26006204";
		wait for Clk_period;
		Addr <=  "0011101101111";
		Trees_din <= x"ff9d1f11";
		wait for Clk_period;
		Addr <=  "0011101110000";
		Trees_din <= x"00541f11";
		wait for Clk_period;
		Addr <=  "0011101110001";
		Trees_din <= x"0800c608";
		wait for Clk_period;
		Addr <=  "0011101110010";
		Trees_din <= x"57fed304";
		wait for Clk_period;
		Addr <=  "0011101110011";
		Trees_din <= x"00121f11";
		wait for Clk_period;
		Addr <=  "0011101110100";
		Trees_din <= x"ffa41f11";
		wait for Clk_period;
		Addr <=  "0011101110101";
		Trees_din <= x"48ff0704";
		wait for Clk_period;
		Addr <=  "0011101110110";
		Trees_din <= x"ffa61f11";
		wait for Clk_period;
		Addr <=  "0011101110111";
		Trees_din <= x"00911f11";
		wait for Clk_period;
		Addr <=  "0011101111000";
		Trees_din <= x"f3fed020";
		wait for Clk_period;
		Addr <=  "0011101111001";
		Trees_din <= x"45ff4f10";
		wait for Clk_period;
		Addr <=  "0011101111010";
		Trees_din <= x"04ffde08";
		wait for Clk_period;
		Addr <=  "0011101111011";
		Trees_din <= x"b1ff6904";
		wait for Clk_period;
		Addr <=  "0011101111100";
		Trees_din <= x"ffa71f11";
		wait for Clk_period;
		Addr <=  "0011101111101";
		Trees_din <= x"004e1f11";
		wait for Clk_period;
		Addr <=  "0011101111110";
		Trees_din <= x"84ffe604";
		wait for Clk_period;
		Addr <=  "0011101111111";
		Trees_din <= x"004d1f11";
		wait for Clk_period;
		Addr <=  "0011110000000";
		Trees_din <= x"000a1f11";
		wait for Clk_period;
		Addr <=  "0011110000001";
		Trees_din <= x"52ff3c08";
		wait for Clk_period;
		Addr <=  "0011110000010";
		Trees_din <= x"7bff2e04";
		wait for Clk_period;
		Addr <=  "0011110000011";
		Trees_din <= x"ffce1f11";
		wait for Clk_period;
		Addr <=  "0011110000100";
		Trees_din <= x"006d1f11";
		wait for Clk_period;
		Addr <=  "0011110000101";
		Trees_din <= x"d6ffbd04";
		wait for Clk_period;
		Addr <=  "0011110000110";
		Trees_din <= x"008f1f11";
		wait for Clk_period;
		Addr <=  "0011110000111";
		Trees_din <= x"ff7a1f11";
		wait for Clk_period;
		Addr <=  "0011110001000";
		Trees_din <= x"26000810";
		wait for Clk_period;
		Addr <=  "0011110001001";
		Trees_din <= x"82ff3d08";
		wait for Clk_period;
		Addr <=  "0011110001010";
		Trees_din <= x"6bff1f04";
		wait for Clk_period;
		Addr <=  "0011110001011";
		Trees_din <= x"00301f11";
		wait for Clk_period;
		Addr <=  "0011110001100";
		Trees_din <= x"ff751f11";
		wait for Clk_period;
		Addr <=  "0011110001101";
		Trees_din <= x"6a002304";
		wait for Clk_period;
		Addr <=  "0011110001110";
		Trees_din <= x"ff6b1f11";
		wait for Clk_period;
		Addr <=  "0011110001111";
		Trees_din <= x"00321f11";
		wait for Clk_period;
		Addr <=  "0011110010000";
		Trees_din <= x"faffc608";
		wait for Clk_period;
		Addr <=  "0011110010001";
		Trees_din <= x"eaff4204";
		wait for Clk_period;
		Addr <=  "0011110010010";
		Trees_din <= x"002a1f11";
		wait for Clk_period;
		Addr <=  "0011110010011";
		Trees_din <= x"ffe01f11";
		wait for Clk_period;
		Addr <=  "0011110010100";
		Trees_din <= x"53feea04";
		wait for Clk_period;
		Addr <=  "0011110010101";
		Trees_din <= x"ff7f1f11";
		wait for Clk_period;
		Addr <=  "0011110010110";
		Trees_din <= x"004f1f11";
		wait for Clk_period;
		Addr <=  "0011110010111";
		Trees_din <= x"d800593c";
		wait for Clk_period;
		Addr <=  "0011110011000";
		Trees_din <= x"09ffcd20";
		wait for Clk_period;
		Addr <=  "0011110011001";
		Trees_din <= x"ddfed810";
		wait for Clk_period;
		Addr <=  "0011110011010";
		Trees_din <= x"baffa208";
		wait for Clk_period;
		Addr <=  "0011110011011";
		Trees_din <= x"f3ff1504";
		wait for Clk_period;
		Addr <=  "0011110011100";
		Trees_din <= x"ff961f11";
		wait for Clk_period;
		Addr <=  "0011110011101";
		Trees_din <= x"00151f11";
		wait for Clk_period;
		Addr <=  "0011110011110";
		Trees_din <= x"75fff604";
		wait for Clk_period;
		Addr <=  "0011110011111";
		Trees_din <= x"fff91f11";
		wait for Clk_period;
		Addr <=  "0011110100000";
		Trees_din <= x"00b31f11";
		wait for Clk_period;
		Addr <=  "0011110100001";
		Trees_din <= x"82ff1208";
		wait for Clk_period;
		Addr <=  "0011110100010";
		Trees_din <= x"17fff504";
		wait for Clk_period;
		Addr <=  "0011110100011";
		Trees_din <= x"008e1f11";
		wait for Clk_period;
		Addr <=  "0011110100100";
		Trees_din <= x"ffa01f11";
		wait for Clk_period;
		Addr <=  "0011110100101";
		Trees_din <= x"65000204";
		wait for Clk_period;
		Addr <=  "0011110100110";
		Trees_din <= x"ff651f11";
		wait for Clk_period;
		Addr <=  "0011110100111";
		Trees_din <= x"00231f11";
		wait for Clk_period;
		Addr <=  "0011110101000";
		Trees_din <= x"4fff3410";
		wait for Clk_period;
		Addr <=  "0011110101001";
		Trees_din <= x"a2ffbe08";
		wait for Clk_period;
		Addr <=  "0011110101010";
		Trees_din <= x"3eff1d04";
		wait for Clk_period;
		Addr <=  "0011110101011";
		Trees_din <= x"fffc1f11";
		wait for Clk_period;
		Addr <=  "0011110101100";
		Trees_din <= x"ff6c1f11";
		wait for Clk_period;
		Addr <=  "0011110101101";
		Trees_din <= x"04002504";
		wait for Clk_period;
		Addr <=  "0011110101110";
		Trees_din <= x"ff9f1f11";
		wait for Clk_period;
		Addr <=  "0011110101111";
		Trees_din <= x"00821f11";
		wait for Clk_period;
		Addr <=  "0011110110000";
		Trees_din <= x"f5005108";
		wait for Clk_period;
		Addr <=  "0011110110001";
		Trees_din <= x"2aff4a04";
		wait for Clk_period;
		Addr <=  "0011110110010";
		Trees_din <= x"ff981f11";
		wait for Clk_period;
		Addr <=  "0011110110011";
		Trees_din <= x"007a1f11";
		wait for Clk_period;
		Addr <=  "0011110110100";
		Trees_din <= x"ff901f11";
		wait for Clk_period;
		Addr <=  "0011110110101";
		Trees_din <= x"c5ff7f14";
		wait for Clk_period;
		Addr <=  "0011110110110";
		Trees_din <= x"8800670c";
		wait for Clk_period;
		Addr <=  "0011110110111";
		Trees_din <= x"f7fe9404";
		wait for Clk_period;
		Addr <=  "0011110111000";
		Trees_din <= x"ffcd1f11";
		wait for Clk_period;
		Addr <=  "0011110111001";
		Trees_din <= x"96ffc004";
		wait for Clk_period;
		Addr <=  "0011110111010";
		Trees_din <= x"00b31f11";
		wait for Clk_period;
		Addr <=  "0011110111011";
		Trees_din <= x"ffed1f11";
		wait for Clk_period;
		Addr <=  "0011110111100";
		Trees_din <= x"62feb704";
		wait for Clk_period;
		Addr <=  "0011110111101";
		Trees_din <= x"00501f11";
		wait for Clk_period;
		Addr <=  "0011110111110";
		Trees_din <= x"ff871f11";
		wait for Clk_period;
		Addr <=  "0011110111111";
		Trees_din <= x"cafe6a04";
		wait for Clk_period;
		Addr <=  "0011111000000";
		Trees_din <= x"ff7f1f11";
		wait for Clk_period;
		Addr <=  "0011111000001";
		Trees_din <= x"83ffc704";
		wait for Clk_period;
		Addr <=  "0011111000010";
		Trees_din <= x"00701f11";
		wait for Clk_period;
		Addr <=  "0011111000011";
		Trees_din <= x"fffa1f11";
		wait for Clk_period;
		Addr <=  "0011111000100";
		Trees_din <= x"60ffbe7c";
		wait for Clk_period;
		Addr <=  "0011111000101";
		Trees_din <= x"3eff8140";
		wait for Clk_period;
		Addr <=  "0011111000110";
		Trees_din <= x"44005320";
		wait for Clk_period;
		Addr <=  "0011111000111";
		Trees_din <= x"3dffe710";
		wait for Clk_period;
		Addr <=  "0011111001000";
		Trees_din <= x"5fff9608";
		wait for Clk_period;
		Addr <=  "0011111001001";
		Trees_din <= x"4efe7f04";
		wait for Clk_period;
		Addr <=  "0011111001010";
		Trees_din <= x"007320c5";
		wait for Clk_period;
		Addr <=  "0011111001011";
		Trees_din <= x"000020c5";
		wait for Clk_period;
		Addr <=  "0011111001100";
		Trees_din <= x"3bff9c04";
		wait for Clk_period;
		Addr <=  "0011111001101";
		Trees_din <= x"ff8920c5";
		wait for Clk_period;
		Addr <=  "0011111001110";
		Trees_din <= x"001d20c5";
		wait for Clk_period;
		Addr <=  "0011111001111";
		Trees_din <= x"f1ff4908";
		wait for Clk_period;
		Addr <=  "0011111010000";
		Trees_din <= x"bf001204";
		wait for Clk_period;
		Addr <=  "0011111010001";
		Trees_din <= x"fffe20c5";
		wait for Clk_period;
		Addr <=  "0011111010010";
		Trees_din <= x"00cd20c5";
		wait for Clk_period;
		Addr <=  "0011111010011";
		Trees_din <= x"19ff3704";
		wait for Clk_period;
		Addr <=  "0011111010100";
		Trees_din <= x"ffef20c5";
		wait for Clk_period;
		Addr <=  "0011111010101";
		Trees_din <= x"ffa620c5";
		wait for Clk_period;
		Addr <=  "0011111010110";
		Trees_din <= x"4eff7d10";
		wait for Clk_period;
		Addr <=  "0011111010111";
		Trees_din <= x"b5feb708";
		wait for Clk_period;
		Addr <=  "0011111011000";
		Trees_din <= x"0bffb304";
		wait for Clk_period;
		Addr <=  "0011111011001";
		Trees_din <= x"ff7820c5";
		wait for Clk_period;
		Addr <=  "0011111011010";
		Trees_din <= x"001a20c5";
		wait for Clk_period;
		Addr <=  "0011111011011";
		Trees_din <= x"29fef804";
		wait for Clk_period;
		Addr <=  "0011111011100";
		Trees_din <= x"ffa120c5";
		wait for Clk_period;
		Addr <=  "0011111011101";
		Trees_din <= x"008220c5";
		wait for Clk_period;
		Addr <=  "0011111011110";
		Trees_din <= x"20ffb208";
		wait for Clk_period;
		Addr <=  "0011111011111";
		Trees_din <= x"71ff8904";
		wait for Clk_period;
		Addr <=  "0011111100000";
		Trees_din <= x"ff8c20c5";
		wait for Clk_period;
		Addr <=  "0011111100001";
		Trees_din <= x"004920c5";
		wait for Clk_period;
		Addr <=  "0011111100010";
		Trees_din <= x"98ff1904";
		wait for Clk_period;
		Addr <=  "0011111100011";
		Trees_din <= x"003920c5";
		wait for Clk_period;
		Addr <=  "0011111100100";
		Trees_din <= x"ff7220c5";
		wait for Clk_period;
		Addr <=  "0011111100101";
		Trees_din <= x"92ff5720";
		wait for Clk_period;
		Addr <=  "0011111100110";
		Trees_din <= x"59ff0d10";
		wait for Clk_period;
		Addr <=  "0011111100111";
		Trees_din <= x"8c007708";
		wait for Clk_period;
		Addr <=  "0011111101000";
		Trees_din <= x"a5fec404";
		wait for Clk_period;
		Addr <=  "0011111101001";
		Trees_din <= x"005620c5";
		wait for Clk_period;
		Addr <=  "0011111101010";
		Trees_din <= x"ff8d20c5";
		wait for Clk_period;
		Addr <=  "0011111101011";
		Trees_din <= x"e3fef704";
		wait for Clk_period;
		Addr <=  "0011111101100";
		Trees_din <= x"006920c5";
		wait for Clk_period;
		Addr <=  "0011111101101";
		Trees_din <= x"ff8620c5";
		wait for Clk_period;
		Addr <=  "0011111101110";
		Trees_din <= x"9bff3d08";
		wait for Clk_period;
		Addr <=  "0011111101111";
		Trees_din <= x"97fed004";
		wait for Clk_period;
		Addr <=  "0011111110000";
		Trees_din <= x"000c20c5";
		wait for Clk_period;
		Addr <=  "0011111110001";
		Trees_din <= x"006e20c5";
		wait for Clk_period;
		Addr <=  "0011111110010";
		Trees_din <= x"81ffd104";
		wait for Clk_period;
		Addr <=  "0011111110011";
		Trees_din <= x"003420c5";
		wait for Clk_period;
		Addr <=  "0011111110100";
		Trees_din <= x"ffcf20c5";
		wait for Clk_period;
		Addr <=  "0011111110101";
		Trees_din <= x"faff150c";
		wait for Clk_period;
		Addr <=  "0011111110110";
		Trees_din <= x"bcff5708";
		wait for Clk_period;
		Addr <=  "0011111110111";
		Trees_din <= x"68fe3c04";
		wait for Clk_period;
		Addr <=  "0011111111000";
		Trees_din <= x"ff9520c5";
		wait for Clk_period;
		Addr <=  "0011111111001";
		Trees_din <= x"009620c5";
		wait for Clk_period;
		Addr <=  "0011111111010";
		Trees_din <= x"ff9420c5";
		wait for Clk_period;
		Addr <=  "0011111111011";
		Trees_din <= x"24ff5a08";
		wait for Clk_period;
		Addr <=  "0011111111100";
		Trees_din <= x"47002504";
		wait for Clk_period;
		Addr <=  "0011111111101";
		Trees_din <= x"ffc520c5";
		wait for Clk_period;
		Addr <=  "0011111111110";
		Trees_din <= x"006e20c5";
		wait for Clk_period;
		Addr <=  "0011111111111";
		Trees_din <= x"01ff8404";
		wait for Clk_period;
		Addr <=  "0100000000000";
		Trees_din <= x"ff8920c5";
		wait for Clk_period;
		Addr <=  "0100000000001";
		Trees_din <= x"008020c5";
		wait for Clk_period;
		Addr <=  "0100000000010";
		Trees_din <= x"05000120";
		wait for Clk_period;
		Addr <=  "0100000000011";
		Trees_din <= x"48000018";
		wait for Clk_period;
		Addr <=  "0100000000100";
		Trees_din <= x"80ff8408";
		wait for Clk_period;
		Addr <=  "0100000000101";
		Trees_din <= x"4dfdfa04";
		wait for Clk_period;
		Addr <=  "0100000000110";
		Trees_din <= x"004320c5";
		wait for Clk_period;
		Addr <=  "0100000000111";
		Trees_din <= x"ff6f20c5";
		wait for Clk_period;
		Addr <=  "0100000001000";
		Trees_din <= x"0dff8f08";
		wait for Clk_period;
		Addr <=  "0100000001001";
		Trees_din <= x"92ff2104";
		wait for Clk_period;
		Addr <=  "0100000001010";
		Trees_din <= x"009120c5";
		wait for Clk_period;
		Addr <=  "0100000001011";
		Trees_din <= x"ffe120c5";
		wait for Clk_period;
		Addr <=  "0100000001100";
		Trees_din <= x"83ff5204";
		wait for Clk_period;
		Addr <=  "0100000001101";
		Trees_din <= x"ff9520c5";
		wait for Clk_period;
		Addr <=  "0100000001110";
		Trees_din <= x"000720c5";
		wait for Clk_period;
		Addr <=  "0100000001111";
		Trees_din <= x"79ffbf04";
		wait for Clk_period;
		Addr <=  "0100000010000";
		Trees_din <= x"ff6820c5";
		wait for Clk_period;
		Addr <=  "0100000010001";
		Trees_din <= x"fffa20c5";
		wait for Clk_period;
		Addr <=  "0100000010010";
		Trees_din <= x"17000320";
		wait for Clk_period;
		Addr <=  "0100000010011";
		Trees_din <= x"7affcc10";
		wait for Clk_period;
		Addr <=  "0100000010100";
		Trees_din <= x"4afeb108";
		wait for Clk_period;
		Addr <=  "0100000010101";
		Trees_din <= x"5eff9e04";
		wait for Clk_period;
		Addr <=  "0100000010110";
		Trees_din <= x"003020c5";
		wait for Clk_period;
		Addr <=  "0100000010111";
		Trees_din <= x"ff7120c5";
		wait for Clk_period;
		Addr <=  "0100000011000";
		Trees_din <= x"94ffcf04";
		wait for Clk_period;
		Addr <=  "0100000011001";
		Trees_din <= x"006420c5";
		wait for Clk_period;
		Addr <=  "0100000011010";
		Trees_din <= x"000620c5";
		wait for Clk_period;
		Addr <=  "0100000011011";
		Trees_din <= x"dfff2a08";
		wait for Clk_period;
		Addr <=  "0100000011100";
		Trees_din <= x"91ffb704";
		wait for Clk_period;
		Addr <=  "0100000011101";
		Trees_din <= x"005920c5";
		wait for Clk_period;
		Addr <=  "0100000011110";
		Trees_din <= x"ffa620c5";
		wait for Clk_period;
		Addr <=  "0100000011111";
		Trees_din <= x"91000004";
		wait for Clk_period;
		Addr <=  "0100000100000";
		Trees_din <= x"00c020c5";
		wait for Clk_period;
		Addr <=  "0100000100001";
		Trees_din <= x"ffe920c5";
		wait for Clk_period;
		Addr <=  "0100000100010";
		Trees_din <= x"73002710";
		wait for Clk_period;
		Addr <=  "0100000100011";
		Trees_din <= x"3bff2e08";
		wait for Clk_period;
		Addr <=  "0100000100100";
		Trees_din <= x"6ffee704";
		wait for Clk_period;
		Addr <=  "0100000100101";
		Trees_din <= x"004920c5";
		wait for Clk_period;
		Addr <=  "0100000100110";
		Trees_din <= x"ff9f20c5";
		wait for Clk_period;
		Addr <=  "0100000100111";
		Trees_din <= x"4eff1e04";
		wait for Clk_period;
		Addr <=  "0100000101000";
		Trees_din <= x"fff320c5";
		wait for Clk_period;
		Addr <=  "0100000101001";
		Trees_din <= x"006620c5";
		wait for Clk_period;
		Addr <=  "0100000101010";
		Trees_din <= x"0a005208";
		wait for Clk_period;
		Addr <=  "0100000101011";
		Trees_din <= x"99ff5c04";
		wait for Clk_period;
		Addr <=  "0100000101100";
		Trees_din <= x"ff5720c5";
		wait for Clk_period;
		Addr <=  "0100000101101";
		Trees_din <= x"002f20c5";
		wait for Clk_period;
		Addr <=  "0100000101110";
		Trees_din <= x"7cff4704";
		wait for Clk_period;
		Addr <=  "0100000101111";
		Trees_din <= x"008a20c5";
		wait for Clk_period;
		Addr <=  "0100000110000";
		Trees_din <= x"ffdf20c5";
		wait for Clk_period;
		Addr <=  "0100000110001";
		Trees_din <= x"6d007068";
		wait for Clk_period;
		Addr <=  "0100000110010";
		Trees_din <= x"6f003e40";
		wait for Clk_period;
		Addr <=  "0100000110011";
		Trees_din <= x"72005220";
		wait for Clk_period;
		Addr <=  "0100000110100";
		Trees_din <= x"8bffb110";
		wait for Clk_period;
		Addr <=  "0100000110101";
		Trees_din <= x"77ff6308";
		wait for Clk_period;
		Addr <=  "0100000110110";
		Trees_din <= x"32ff7904";
		wait for Clk_period;
		Addr <=  "0100000110111";
		Trees_din <= x"006921e1";
		wait for Clk_period;
		Addr <=  "0100000111000";
		Trees_din <= x"ffd321e1";
		wait for Clk_period;
		Addr <=  "0100000111001";
		Trees_din <= x"adffc104";
		wait for Clk_period;
		Addr <=  "0100000111010";
		Trees_din <= x"ff7b21e1";
		wait for Clk_period;
		Addr <=  "0100000111011";
		Trees_din <= x"003521e1";
		wait for Clk_period;
		Addr <=  "0100000111100";
		Trees_din <= x"b1ff2a08";
		wait for Clk_period;
		Addr <=  "0100000111101";
		Trees_din <= x"86fef304";
		wait for Clk_period;
		Addr <=  "0100000111110";
		Trees_din <= x"fff721e1";
		wait for Clk_period;
		Addr <=  "0100000111111";
		Trees_din <= x"ffbd21e1";
		wait for Clk_period;
		Addr <=  "0100001000000";
		Trees_din <= x"b4ff6104";
		wait for Clk_period;
		Addr <=  "0100001000001";
		Trees_din <= x"001a21e1";
		wait for Clk_period;
		Addr <=  "0100001000010";
		Trees_din <= x"ffcd21e1";
		wait for Clk_period;
		Addr <=  "0100001000011";
		Trees_din <= x"74fffc10";
		wait for Clk_period;
		Addr <=  "0100001000100";
		Trees_din <= x"29ff8108";
		wait for Clk_period;
		Addr <=  "0100001000101";
		Trees_din <= x"5bffa604";
		wait for Clk_period;
		Addr <=  "0100001000110";
		Trees_din <= x"007421e1";
		wait for Clk_period;
		Addr <=  "0100001000111";
		Trees_din <= x"ffdd21e1";
		wait for Clk_period;
		Addr <=  "0100001001000";
		Trees_din <= x"e9fee804";
		wait for Clk_period;
		Addr <=  "0100001001001";
		Trees_din <= x"003721e1";
		wait for Clk_period;
		Addr <=  "0100001001010";
		Trees_din <= x"ffd421e1";
		wait for Clk_period;
		Addr <=  "0100001001011";
		Trees_din <= x"22011c08";
		wait for Clk_period;
		Addr <=  "0100001001100";
		Trees_din <= x"49005504";
		wait for Clk_period;
		Addr <=  "0100001001101";
		Trees_din <= x"ffbe21e1";
		wait for Clk_period;
		Addr <=  "0100001001110";
		Trees_din <= x"003a21e1";
		wait for Clk_period;
		Addr <=  "0100001001111";
		Trees_din <= x"cbffda04";
		wait for Clk_period;
		Addr <=  "0100001010000";
		Trees_din <= x"009321e1";
		wait for Clk_period;
		Addr <=  "0100001010001";
		Trees_din <= x"ffce21e1";
		wait for Clk_period;
		Addr <=  "0100001010010";
		Trees_din <= x"15ffb918";
		wait for Clk_period;
		Addr <=  "0100001010011";
		Trees_din <= x"29ffba10";
		wait for Clk_period;
		Addr <=  "0100001010100";
		Trees_din <= x"9eff6008";
		wait for Clk_period;
		Addr <=  "0100001010101";
		Trees_din <= x"31ffa604";
		wait for Clk_period;
		Addr <=  "0100001010110";
		Trees_din <= x"ffaa21e1";
		wait for Clk_period;
		Addr <=  "0100001010111";
		Trees_din <= x"006f21e1";
		wait for Clk_period;
		Addr <=  "0100001011000";
		Trees_din <= x"a5feb404";
		wait for Clk_period;
		Addr <=  "0100001011001";
		Trees_din <= x"ffe221e1";
		wait for Clk_period;
		Addr <=  "0100001011010";
		Trees_din <= x"00a521e1";
		wait for Clk_period;
		Addr <=  "0100001011011";
		Trees_din <= x"92ff3304";
		wait for Clk_period;
		Addr <=  "0100001011100";
		Trees_din <= x"ff9a21e1";
		wait for Clk_period;
		Addr <=  "0100001011101";
		Trees_din <= x"000f21e1";
		wait for Clk_period;
		Addr <=  "0100001011110";
		Trees_din <= x"8ffec908";
		wait for Clk_period;
		Addr <=  "0100001011111";
		Trees_din <= x"82ff4404";
		wait for Clk_period;
		Addr <=  "0100001100000";
		Trees_din <= x"ffde21e1";
		wait for Clk_period;
		Addr <=  "0100001100001";
		Trees_din <= x"ff7a21e1";
		wait for Clk_period;
		Addr <=  "0100001100010";
		Trees_din <= x"75002a04";
		wait for Clk_period;
		Addr <=  "0100001100011";
		Trees_din <= x"007021e1";
		wait for Clk_period;
		Addr <=  "0100001100100";
		Trees_din <= x"fffd21e1";
		wait for Clk_period;
		Addr <=  "0100001100101";
		Trees_din <= x"20ff1510";
		wait for Clk_period;
		Addr <=  "0100001100110";
		Trees_din <= x"cafe0608";
		wait for Clk_period;
		Addr <=  "0100001100111";
		Trees_din <= x"a0ff3604";
		wait for Clk_period;
		Addr <=  "0100001101000";
		Trees_din <= x"ffc221e1";
		wait for Clk_period;
		Addr <=  "0100001101001";
		Trees_din <= x"008121e1";
		wait for Clk_period;
		Addr <=  "0100001101010";
		Trees_din <= x"a9000604";
		wait for Clk_period;
		Addr <=  "0100001101011";
		Trees_din <= x"ff6b21e1";
		wait for Clk_period;
		Addr <=  "0100001101100";
		Trees_din <= x"003c21e1";
		wait for Clk_period;
		Addr <=  "0100001101101";
		Trees_din <= x"f1006f14";
		wait for Clk_period;
		Addr <=  "0100001101110";
		Trees_din <= x"50fe2b04";
		wait for Clk_period;
		Addr <=  "0100001101111";
		Trees_din <= x"ff7f21e1";
		wait for Clk_period;
		Addr <=  "0100001110000";
		Trees_din <= x"4dfdaf08";
		wait for Clk_period;
		Addr <=  "0100001110001";
		Trees_din <= x"1dff0004";
		wait for Clk_period;
		Addr <=  "0100001110010";
		Trees_din <= x"ff7c21e1";
		wait for Clk_period;
		Addr <=  "0100001110011";
		Trees_din <= x"ffe521e1";
		wait for Clk_period;
		Addr <=  "0100001110100";
		Trees_din <= x"8800ba04";
		wait for Clk_period;
		Addr <=  "0100001110101";
		Trees_din <= x"004721e1";
		wait for Clk_period;
		Addr <=  "0100001110110";
		Trees_din <= x"ffe721e1";
		wait for Clk_period;
		Addr <=  "0100001110111";
		Trees_din <= x"ff8921e1";
		wait for Clk_period;
		Addr <=  "0100001111000";
		Trees_din <= x"33ff5a64";
		wait for Clk_period;
		Addr <=  "0100001111001";
		Trees_din <= x"62ff4530";
		wait for Clk_period;
		Addr <=  "0100001111010";
		Trees_din <= x"77ffbc1c";
		wait for Clk_period;
		Addr <=  "0100001111011";
		Trees_din <= x"e3ff3110";
		wait for Clk_period;
		Addr <=  "0100001111100";
		Trees_din <= x"7afff708";
		wait for Clk_period;
		Addr <=  "0100001111101";
		Trees_din <= x"c2002d04";
		wait for Clk_period;
		Addr <=  "0100001111110";
		Trees_din <= x"002723a5";
		wait for Clk_period;
		Addr <=  "0100001111111";
		Trees_din <= x"ffab23a5";
		wait for Clk_period;
		Addr <=  "0100010000000";
		Trees_din <= x"9eff3c04";
		wait for Clk_period;
		Addr <=  "0100010000001";
		Trees_din <= x"fff723a5";
		wait for Clk_period;
		Addr <=  "0100010000010";
		Trees_din <= x"008d23a5";
		wait for Clk_period;
		Addr <=  "0100010000011";
		Trees_din <= x"bf000208";
		wait for Clk_period;
		Addr <=  "0100010000100";
		Trees_din <= x"41ff5604";
		wait for Clk_period;
		Addr <=  "0100010000101";
		Trees_din <= x"ff6e23a5";
		wait for Clk_period;
		Addr <=  "0100010000110";
		Trees_din <= x"001323a5";
		wait for Clk_period;
		Addr <=  "0100010000111";
		Trees_din <= x"005923a5";
		wait for Clk_period;
		Addr <=  "0100010001000";
		Trees_din <= x"0800eb0c";
		wait for Clk_period;
		Addr <=  "0100010001001";
		Trees_din <= x"d1fee604";
		wait for Clk_period;
		Addr <=  "0100010001010";
		Trees_din <= x"001723a5";
		wait for Clk_period;
		Addr <=  "0100010001011";
		Trees_din <= x"cc001804";
		wait for Clk_period;
		Addr <=  "0100010001100";
		Trees_din <= x"ff6823a5";
		wait for Clk_period;
		Addr <=  "0100010001101";
		Trees_din <= x"fffa23a5";
		wait for Clk_period;
		Addr <=  "0100010001110";
		Trees_din <= x"12003004";
		wait for Clk_period;
		Addr <=  "0100010001111";
		Trees_din <= x"004d23a5";
		wait for Clk_period;
		Addr <=  "0100010010000";
		Trees_din <= x"ffd023a5";
		wait for Clk_period;
		Addr <=  "0100010010001";
		Trees_din <= x"85ff0818";
		wait for Clk_period;
		Addr <=  "0100010010010";
		Trees_din <= x"4fff550c";
		wait for Clk_period;
		Addr <=  "0100010010011";
		Trees_din <= x"a4ff3404";
		wait for Clk_period;
		Addr <=  "0100010010100";
		Trees_din <= x"007823a5";
		wait for Clk_period;
		Addr <=  "0100010010101";
		Trees_din <= x"3bff3004";
		wait for Clk_period;
		Addr <=  "0100010010110";
		Trees_din <= x"fff423a5";
		wait for Clk_period;
		Addr <=  "0100010010111";
		Trees_din <= x"ff7723a5";
		wait for Clk_period;
		Addr <=  "0100010011000";
		Trees_din <= x"e3fe6804";
		wait for Clk_period;
		Addr <=  "0100010011001";
		Trees_din <= x"ffad23a5";
		wait for Clk_period;
		Addr <=  "0100010011010";
		Trees_din <= x"ddfea404";
		wait for Clk_period;
		Addr <=  "0100010011011";
		Trees_din <= x"ffc623a5";
		wait for Clk_period;
		Addr <=  "0100010011100";
		Trees_din <= x"009623a5";
		wait for Clk_period;
		Addr <=  "0100010011101";
		Trees_din <= x"c5ff8b10";
		wait for Clk_period;
		Addr <=  "0100010011110";
		Trees_din <= x"84ffd008";
		wait for Clk_period;
		Addr <=  "0100010011111";
		Trees_din <= x"9dff1904";
		wait for Clk_period;
		Addr <=  "0100010100000";
		Trees_din <= x"005823a5";
		wait for Clk_period;
		Addr <=  "0100010100001";
		Trees_din <= x"fff523a5";
		wait for Clk_period;
		Addr <=  "0100010100010";
		Trees_din <= x"5bff6004";
		wait for Clk_period;
		Addr <=  "0100010100011";
		Trees_din <= x"fff023a5";
		wait for Clk_period;
		Addr <=  "0100010100100";
		Trees_din <= x"ff8723a5";
		wait for Clk_period;
		Addr <=  "0100010100101";
		Trees_din <= x"6d008108";
		wait for Clk_period;
		Addr <=  "0100010100110";
		Trees_din <= x"0cfdf904";
		wait for Clk_period;
		Addr <=  "0100010100111";
		Trees_din <= x"fff823a5";
		wait for Clk_period;
		Addr <=  "0100010101000";
		Trees_din <= x"ff6423a5";
		wait for Clk_period;
		Addr <=  "0100010101001";
		Trees_din <= x"002723a5";
		wait for Clk_period;
		Addr <=  "0100010101010";
		Trees_din <= x"b0ff4f40";
		wait for Clk_period;
		Addr <=  "0100010101011";
		Trees_din <= x"32feea20";
		wait for Clk_period;
		Addr <=  "0100010101100";
		Trees_din <= x"dcffe810";
		wait for Clk_period;
		Addr <=  "0100010101101";
		Trees_din <= x"5dff4f08";
		wait for Clk_period;
		Addr <=  "0100010101110";
		Trees_din <= x"82ff1204";
		wait for Clk_period;
		Addr <=  "0100010101111";
		Trees_din <= x"ff9523a5";
		wait for Clk_period;
		Addr <=  "0100010110000";
		Trees_din <= x"008223a5";
		wait for Clk_period;
		Addr <=  "0100010110001";
		Trees_din <= x"d5ffcd04";
		wait for Clk_period;
		Addr <=  "0100010110010";
		Trees_din <= x"ff6223a5";
		wait for Clk_period;
		Addr <=  "0100010110011";
		Trees_din <= x"ffd823a5";
		wait for Clk_period;
		Addr <=  "0100010110100";
		Trees_din <= x"58ff1e08";
		wait for Clk_period;
		Addr <=  "0100010110101";
		Trees_din <= x"9affa304";
		wait for Clk_period;
		Addr <=  "0100010110110";
		Trees_din <= x"ffae23a5";
		wait for Clk_period;
		Addr <=  "0100010110111";
		Trees_din <= x"007423a5";
		wait for Clk_period;
		Addr <=  "0100010111000";
		Trees_din <= x"98fe5204";
		wait for Clk_period;
		Addr <=  "0100010111001";
		Trees_din <= x"004423a5";
		wait for Clk_period;
		Addr <=  "0100010111010";
		Trees_din <= x"ff8523a5";
		wait for Clk_period;
		Addr <=  "0100010111011";
		Trees_din <= x"55003b10";
		wait for Clk_period;
		Addr <=  "0100010111100";
		Trees_din <= x"47ff3e08";
		wait for Clk_period;
		Addr <=  "0100010111101";
		Trees_din <= x"15ff9504";
		wait for Clk_period;
		Addr <=  "0100010111110";
		Trees_din <= x"ff7c23a5";
		wait for Clk_period;
		Addr <=  "0100010111111";
		Trees_din <= x"001823a5";
		wait for Clk_period;
		Addr <=  "0100011000000";
		Trees_din <= x"3d006404";
		wait for Clk_period;
		Addr <=  "0100011000001";
		Trees_din <= x"007323a5";
		wait for Clk_period;
		Addr <=  "0100011000010";
		Trees_din <= x"ff8b23a5";
		wait for Clk_period;
		Addr <=  "0100011000011";
		Trees_din <= x"27ff9208";
		wait for Clk_period;
		Addr <=  "0100011000100";
		Trees_din <= x"ceff9e04";
		wait for Clk_period;
		Addr <=  "0100011000101";
		Trees_din <= x"ffd623a5";
		wait for Clk_period;
		Addr <=  "0100011000110";
		Trees_din <= x"00c223a5";
		wait for Clk_period;
		Addr <=  "0100011000111";
		Trees_din <= x"af001204";
		wait for Clk_period;
		Addr <=  "0100011001000";
		Trees_din <= x"ff7a23a5";
		wait for Clk_period;
		Addr <=  "0100011001001";
		Trees_din <= x"006623a5";
		wait for Clk_period;
		Addr <=  "0100011001010";
		Trees_din <= x"79fed120";
		wait for Clk_period;
		Addr <=  "0100011001011";
		Trees_din <= x"53ff8310";
		wait for Clk_period;
		Addr <=  "0100011001100";
		Trees_din <= x"4eff0908";
		wait for Clk_period;
		Addr <=  "0100011001101";
		Trees_din <= x"ec001004";
		wait for Clk_period;
		Addr <=  "0100011001110";
		Trees_din <= x"ffb523a5";
		wait for Clk_period;
		Addr <=  "0100011001111";
		Trees_din <= x"008923a5";
		wait for Clk_period;
		Addr <=  "0100011010000";
		Trees_din <= x"b5ff7704";
		wait for Clk_period;
		Addr <=  "0100011010001";
		Trees_din <= x"ff6423a5";
		wait for Clk_period;
		Addr <=  "0100011010010";
		Trees_din <= x"000723a5";
		wait for Clk_period;
		Addr <=  "0100011010011";
		Trees_din <= x"15ff9a08";
		wait for Clk_period;
		Addr <=  "0100011010100";
		Trees_din <= x"26001804";
		wait for Clk_period;
		Addr <=  "0100011010101";
		Trees_din <= x"fff123a5";
		wait for Clk_period;
		Addr <=  "0100011010110";
		Trees_din <= x"00b523a5";
		wait for Clk_period;
		Addr <=  "0100011010111";
		Trees_din <= x"28ff5004";
		wait for Clk_period;
		Addr <=  "0100011011000";
		Trees_din <= x"ff9b23a5";
		wait for Clk_period;
		Addr <=  "0100011011001";
		Trees_din <= x"005d23a5";
		wait for Clk_period;
		Addr <=  "0100011011010";
		Trees_din <= x"2bffd910";
		wait for Clk_period;
		Addr <=  "0100011011011";
		Trees_din <= x"fbffd708";
		wait for Clk_period;
		Addr <=  "0100011011100";
		Trees_din <= x"0cfdbd04";
		wait for Clk_period;
		Addr <=  "0100011011101";
		Trees_din <= x"006e23a5";
		wait for Clk_period;
		Addr <=  "0100011011110";
		Trees_din <= x"ffc123a5";
		wait for Clk_period;
		Addr <=  "0100011011111";
		Trees_din <= x"43ff9b04";
		wait for Clk_period;
		Addr <=  "0100011100000";
		Trees_din <= x"003923a5";
		wait for Clk_period;
		Addr <=  "0100011100001";
		Trees_din <= x"ff9b23a5";
		wait for Clk_period;
		Addr <=  "0100011100010";
		Trees_din <= x"e4ff7e08";
		wait for Clk_period;
		Addr <=  "0100011100011";
		Trees_din <= x"db00e604";
		wait for Clk_period;
		Addr <=  "0100011100100";
		Trees_din <= x"ff8a23a5";
		wait for Clk_period;
		Addr <=  "0100011100101";
		Trees_din <= x"006423a5";
		wait for Clk_period;
		Addr <=  "0100011100110";
		Trees_din <= x"92ff2404";
		wait for Clk_period;
		Addr <=  "0100011100111";
		Trees_din <= x"00ac23a5";
		wait for Clk_period;
		Addr <=  "0100011101000";
		Trees_din <= x"ffa523a5";
		wait for Clk_period;
		Addr <=  "0100011101001";
		Trees_din <= x"2eff5274";
		wait for Clk_period;
		Addr <=  "0100011101010";
		Trees_din <= x"24ffb840";
		wait for Clk_period;
		Addr <=  "0100011101011";
		Trees_din <= x"6fff7520";
		wait for Clk_period;
		Addr <=  "0100011101100";
		Trees_din <= x"2eff4010";
		wait for Clk_period;
		Addr <=  "0100011101101";
		Trees_din <= x"0dff4a08";
		wait for Clk_period;
		Addr <=  "0100011101110";
		Trees_din <= x"b5ff0204";
		wait for Clk_period;
		Addr <=  "0100011101111";
		Trees_din <= x"00662561";
		wait for Clk_period;
		Addr <=  "0100011110000";
		Trees_din <= x"ffd12561";
		wait for Clk_period;
		Addr <=  "0100011110001";
		Trees_din <= x"ebff4504";
		wait for Clk_period;
		Addr <=  "0100011110010";
		Trees_din <= x"ffaa2561";
		wait for Clk_period;
		Addr <=  "0100011110011";
		Trees_din <= x"00592561";
		wait for Clk_period;
		Addr <=  "0100011110100";
		Trees_din <= x"00ff8e08";
		wait for Clk_period;
		Addr <=  "0100011110101";
		Trees_din <= x"b4ff9904";
		wait for Clk_period;
		Addr <=  "0100011110110";
		Trees_din <= x"00942561";
		wait for Clk_period;
		Addr <=  "0100011110111";
		Trees_din <= x"ffef2561";
		wait for Clk_period;
		Addr <=  "0100011111000";
		Trees_din <= x"87ff2a04";
		wait for Clk_period;
		Addr <=  "0100011111001";
		Trees_din <= x"00392561";
		wait for Clk_period;
		Addr <=  "0100011111010";
		Trees_din <= x"ff972561";
		wait for Clk_period;
		Addr <=  "0100011111011";
		Trees_din <= x"aaff8310";
		wait for Clk_period;
		Addr <=  "0100011111100";
		Trees_din <= x"cfffbe08";
		wait for Clk_period;
		Addr <=  "0100011111101";
		Trees_din <= x"7dffb004";
		wait for Clk_period;
		Addr <=  "0100011111110";
		Trees_din <= x"ffb92561";
		wait for Clk_period;
		Addr <=  "0100011111111";
		Trees_din <= x"00612561";
		wait for Clk_period;
		Addr <=  "0100100000000";
		Trees_din <= x"fcfedd04";
		wait for Clk_period;
		Addr <=  "0100100000001";
		Trees_din <= x"ffe42561";
		wait for Clk_period;
		Addr <=  "0100100000010";
		Trees_din <= x"00ad2561";
		wait for Clk_period;
		Addr <=  "0100100000011";
		Trees_din <= x"b0ff3c08";
		wait for Clk_period;
		Addr <=  "0100100000100";
		Trees_din <= x"feffff04";
		wait for Clk_period;
		Addr <=  "0100100000101";
		Trees_din <= x"ff892561";
		wait for Clk_period;
		Addr <=  "0100100000110";
		Trees_din <= x"00292561";
		wait for Clk_period;
		Addr <=  "0100100000111";
		Trees_din <= x"d3ff2e04";
		wait for Clk_period;
		Addr <=  "0100100001000";
		Trees_din <= x"007d2561";
		wait for Clk_period;
		Addr <=  "0100100001001";
		Trees_din <= x"ffd12561";
		wait for Clk_period;
		Addr <=  "0100100001010";
		Trees_din <= x"7fff1318";
		wait for Clk_period;
		Addr <=  "0100100001011";
		Trees_din <= x"bf000c10";
		wait for Clk_period;
		Addr <=  "0100100001100";
		Trees_din <= x"5a00ea08";
		wait for Clk_period;
		Addr <=  "0100100001101";
		Trees_din <= x"93ffe104";
		wait for Clk_period;
		Addr <=  "0100100001110";
		Trees_din <= x"ffa32561";
		wait for Clk_period;
		Addr <=  "0100100001111";
		Trees_din <= x"00522561";
		wait for Clk_period;
		Addr <=  "0100100010000";
		Trees_din <= x"4fff4804";
		wait for Clk_period;
		Addr <=  "0100100010001";
		Trees_din <= x"ffd02561";
		wait for Clk_period;
		Addr <=  "0100100010010";
		Trees_din <= x"009c2561";
		wait for Clk_period;
		Addr <=  "0100100010011";
		Trees_din <= x"c7ff0904";
		wait for Clk_period;
		Addr <=  "0100100010100";
		Trees_din <= x"00ca2561";
		wait for Clk_period;
		Addr <=  "0100100010101";
		Trees_din <= x"00012561";
		wait for Clk_period;
		Addr <=  "0100100010110";
		Trees_din <= x"1cff6610";
		wait for Clk_period;
		Addr <=  "0100100010111";
		Trees_din <= x"6fffaa08";
		wait for Clk_period;
		Addr <=  "0100100011000";
		Trees_din <= x"74ffc404";
		wait for Clk_period;
		Addr <=  "0100100011001";
		Trees_din <= x"003d2561";
		wait for Clk_period;
		Addr <=  "0100100011010";
		Trees_din <= x"ff7a2561";
		wait for Clk_period;
		Addr <=  "0100100011011";
		Trees_din <= x"8cffbf04";
		wait for Clk_period;
		Addr <=  "0100100011100";
		Trees_din <= x"ffbe2561";
		wait for Clk_period;
		Addr <=  "0100100011101";
		Trees_din <= x"00a42561";
		wait for Clk_period;
		Addr <=  "0100100011110";
		Trees_din <= x"46fe7f04";
		wait for Clk_period;
		Addr <=  "0100100011111";
		Trees_din <= x"00672561";
		wait for Clk_period;
		Addr <=  "0100100100000";
		Trees_din <= x"d2ff8804";
		wait for Clk_period;
		Addr <=  "0100100100001";
		Trees_din <= x"ff692561";
		wait for Clk_period;
		Addr <=  "0100100100010";
		Trees_din <= x"00242561";
		wait for Clk_period;
		Addr <=  "0100100100011";
		Trees_din <= x"d700ff40";
		wait for Clk_period;
		Addr <=  "0100100100100";
		Trees_din <= x"25000f20";
		wait for Clk_period;
		Addr <=  "0100100100101";
		Trees_din <= x"31006710";
		wait for Clk_period;
		Addr <=  "0100100100110";
		Trees_din <= x"ddff4e08";
		wait for Clk_period;
		Addr <=  "0100100100111";
		Trees_din <= x"83ffa504";
		wait for Clk_period;
		Addr <=  "0100100101000";
		Trees_din <= x"ffdd2561";
		wait for Clk_period;
		Addr <=  "0100100101001";
		Trees_din <= x"00402561";
		wait for Clk_period;
		Addr <=  "0100100101010";
		Trees_din <= x"7cff1604";
		wait for Clk_period;
		Addr <=  "0100100101011";
		Trees_din <= x"00442561";
		wait for Clk_period;
		Addr <=  "0100100101100";
		Trees_din <= x"ff9c2561";
		wait for Clk_period;
		Addr <=  "0100100101101";
		Trees_din <= x"f4fe8708";
		wait for Clk_period;
		Addr <=  "0100100101110";
		Trees_din <= x"ebfea104";
		wait for Clk_period;
		Addr <=  "0100100101111";
		Trees_din <= x"003b2561";
		wait for Clk_period;
		Addr <=  "0100100110000";
		Trees_din <= x"ff722561";
		wait for Clk_period;
		Addr <=  "0100100110001";
		Trees_din <= x"34fff204";
		wait for Clk_period;
		Addr <=  "0100100110010";
		Trees_din <= x"ffd12561";
		wait for Clk_period;
		Addr <=  "0100100110011";
		Trees_din <= x"00612561";
		wait for Clk_period;
		Addr <=  "0100100110100";
		Trees_din <= x"45ff2510";
		wait for Clk_period;
		Addr <=  "0100100110101";
		Trees_din <= x"dc004608";
		wait for Clk_period;
		Addr <=  "0100100110110";
		Trees_din <= x"21006a04";
		wait for Clk_period;
		Addr <=  "0100100110111";
		Trees_din <= x"00212561";
		wait for Clk_period;
		Addr <=  "0100100111000";
		Trees_din <= x"ff882561";
		wait for Clk_period;
		Addr <=  "0100100111001";
		Trees_din <= x"aefee204";
		wait for Clk_period;
		Addr <=  "0100100111010";
		Trees_din <= x"00142561";
		wait for Clk_period;
		Addr <=  "0100100111011";
		Trees_din <= x"ffad2561";
		wait for Clk_period;
		Addr <=  "0100100111100";
		Trees_din <= x"36fff908";
		wait for Clk_period;
		Addr <=  "0100100111101";
		Trees_din <= x"63ffa404";
		wait for Clk_period;
		Addr <=  "0100100111110";
		Trees_din <= x"ffb12561";
		wait for Clk_period;
		Addr <=  "0100100111111";
		Trees_din <= x"000f2561";
		wait for Clk_period;
		Addr <=  "0100101000000";
		Trees_din <= x"80ffca04";
		wait for Clk_period;
		Addr <=  "0100101000001";
		Trees_din <= x"00852561";
		wait for Clk_period;
		Addr <=  "0100101000010";
		Trees_din <= x"ff892561";
		wait for Clk_period;
		Addr <=  "0100101000011";
		Trees_din <= x"b6ff4914";
		wait for Clk_period;
		Addr <=  "0100101000100";
		Trees_din <= x"d600d80c";
		wait for Clk_period;
		Addr <=  "0100101000101";
		Trees_din <= x"6bff0308";
		wait for Clk_period;
		Addr <=  "0100101000110";
		Trees_din <= x"bdff1b04";
		wait for Clk_period;
		Addr <=  "0100101000111";
		Trees_din <= x"00002561";
		wait for Clk_period;
		Addr <=  "0100101001000";
		Trees_din <= x"ff642561";
		wait for Clk_period;
		Addr <=  "0100101001001";
		Trees_din <= x"006b2561";
		wait for Clk_period;
		Addr <=  "0100101001010";
		Trees_din <= x"1dff2404";
		wait for Clk_period;
		Addr <=  "0100101001011";
		Trees_din <= x"00162561";
		wait for Clk_period;
		Addr <=  "0100101001100";
		Trees_din <= x"007f2561";
		wait for Clk_period;
		Addr <=  "0100101001101";
		Trees_din <= x"02fe3c08";
		wait for Clk_period;
		Addr <=  "0100101001110";
		Trees_din <= x"bcfec504";
		wait for Clk_period;
		Addr <=  "0100101001111";
		Trees_din <= x"00362561";
		wait for Clk_period;
		Addr <=  "0100101010000";
		Trees_din <= x"ff902561";
		wait for Clk_period;
		Addr <=  "0100101010001";
		Trees_din <= x"53ff6208";
		wait for Clk_period;
		Addr <=  "0100101010010";
		Trees_din <= x"ab005704";
		wait for Clk_period;
		Addr <=  "0100101010011";
		Trees_din <= x"00512561";
		wait for Clk_period;
		Addr <=  "0100101010100";
		Trees_din <= x"ff942561";
		wait for Clk_period;
		Addr <=  "0100101010101";
		Trees_din <= x"49ff9a04";
		wait for Clk_period;
		Addr <=  "0100101010110";
		Trees_din <= x"ffc02561";
		wait for Clk_period;
		Addr <=  "0100101010111";
		Trees_din <= x"00a02561";
		wait for Clk_period;
		Addr <=  "0100101011000";
		Trees_din <= x"55008374";
		wait for Clk_period;
		Addr <=  "0100101011001";
		Trees_din <= x"a0ff6540";
		wait for Clk_period;
		Addr <=  "0100101011010";
		Trees_din <= x"5dffe120";
		wait for Clk_period;
		Addr <=  "0100101011011";
		Trees_din <= x"b7ff3a10";
		wait for Clk_period;
		Addr <=  "0100101011100";
		Trees_din <= x"c3000f08";
		wait for Clk_period;
		Addr <=  "0100101011101";
		Trees_din <= x"20001d04";
		wait for Clk_period;
		Addr <=  "0100101011110";
		Trees_din <= x"ff9a26fd";
		wait for Clk_period;
		Addr <=  "0100101011111";
		Trees_din <= x"001a26fd";
		wait for Clk_period;
		Addr <=  "0100101100000";
		Trees_din <= x"7dffa004";
		wait for Clk_period;
		Addr <=  "0100101100001";
		Trees_din <= x"ff8f26fd";
		wait for Clk_period;
		Addr <=  "0100101100010";
		Trees_din <= x"004626fd";
		wait for Clk_period;
		Addr <=  "0100101100011";
		Trees_din <= x"d3ff5208";
		wait for Clk_period;
		Addr <=  "0100101100100";
		Trees_din <= x"9cfeb604";
		wait for Clk_period;
		Addr <=  "0100101100101";
		Trees_din <= x"006926fd";
		wait for Clk_period;
		Addr <=  "0100101100110";
		Trees_din <= x"000f26fd";
		wait for Clk_period;
		Addr <=  "0100101100111";
		Trees_din <= x"0aff9f04";
		wait for Clk_period;
		Addr <=  "0100101101000";
		Trees_din <= x"ffe726fd";
		wait for Clk_period;
		Addr <=  "0100101101001";
		Trees_din <= x"006026fd";
		wait for Clk_period;
		Addr <=  "0100101101010";
		Trees_din <= x"6bfea610";
		wait for Clk_period;
		Addr <=  "0100101101011";
		Trees_din <= x"95ff1f08";
		wait for Clk_period;
		Addr <=  "0100101101100";
		Trees_din <= x"d3febe04";
		wait for Clk_period;
		Addr <=  "0100101101101";
		Trees_din <= x"ffe626fd";
		wait for Clk_period;
		Addr <=  "0100101101110";
		Trees_din <= x"005c26fd";
		wait for Clk_period;
		Addr <=  "0100101101111";
		Trees_din <= x"a4ff4504";
		wait for Clk_period;
		Addr <=  "0100101110000";
		Trees_din <= x"005d26fd";
		wait for Clk_period;
		Addr <=  "0100101110001";
		Trees_din <= x"ffb226fd";
		wait for Clk_period;
		Addr <=  "0100101110010";
		Trees_din <= x"afff4208";
		wait for Clk_period;
		Addr <=  "0100101110011";
		Trees_din <= x"59000004";
		wait for Clk_period;
		Addr <=  "0100101110100";
		Trees_din <= x"fff626fd";
		wait for Clk_period;
		Addr <=  "0100101110101";
		Trees_din <= x"007926fd";
		wait for Clk_period;
		Addr <=  "0100101110110";
		Trees_din <= x"0bff0e04";
		wait for Clk_period;
		Addr <=  "0100101110111";
		Trees_din <= x"006426fd";
		wait for Clk_period;
		Addr <=  "0100101111000";
		Trees_din <= x"ffbe26fd";
		wait for Clk_period;
		Addr <=  "0100101111001";
		Trees_din <= x"81ff4f18";
		wait for Clk_period;
		Addr <=  "0100101111010";
		Trees_din <= x"97ff3a10";
		wait for Clk_period;
		Addr <=  "0100101111011";
		Trees_din <= x"0400bb08";
		wait for Clk_period;
		Addr <=  "0100101111100";
		Trees_din <= x"4bfe9f04";
		wait for Clk_period;
		Addr <=  "0100101111101";
		Trees_din <= x"002726fd";
		wait for Clk_period;
		Addr <=  "0100101111110";
		Trees_din <= x"ff8926fd";
		wait for Clk_period;
		Addr <=  "0100101111111";
		Trees_din <= x"54008c04";
		wait for Clk_period;
		Addr <=  "0100110000000";
		Trees_din <= x"001626fd";
		wait for Clk_period;
		Addr <=  "0100110000001";
		Trees_din <= x"005d26fd";
		wait for Clk_period;
		Addr <=  "0100110000010";
		Trees_din <= x"bdffe504";
		wait for Clk_period;
		Addr <=  "0100110000011";
		Trees_din <= x"009026fd";
		wait for Clk_period;
		Addr <=  "0100110000100";
		Trees_din <= x"ffdc26fd";
		wait for Clk_period;
		Addr <=  "0100110000101";
		Trees_din <= x"0fffe510";
		wait for Clk_period;
		Addr <=  "0100110000110";
		Trees_din <= x"6f002c08";
		wait for Clk_period;
		Addr <=  "0100110000111";
		Trees_din <= x"08013804";
		wait for Clk_period;
		Addr <=  "0100110001000";
		Trees_din <= x"ff9b26fd";
		wait for Clk_period;
		Addr <=  "0100110001001";
		Trees_din <= x"005e26fd";
		wait for Clk_period;
		Addr <=  "0100110001010";
		Trees_din <= x"acffcd04";
		wait for Clk_period;
		Addr <=  "0100110001011";
		Trees_din <= x"007926fd";
		wait for Clk_period;
		Addr <=  "0100110001100";
		Trees_din <= x"fff426fd";
		wait for Clk_period;
		Addr <=  "0100110001101";
		Trees_din <= x"f5001808";
		wait for Clk_period;
		Addr <=  "0100110001110";
		Trees_din <= x"14ff1604";
		wait for Clk_period;
		Addr <=  "0100110001111";
		Trees_din <= x"ffd126fd";
		wait for Clk_period;
		Addr <=  "0100110010000";
		Trees_din <= x"007e26fd";
		wait for Clk_period;
		Addr <=  "0100110010001";
		Trees_din <= x"ffaa26fd";
		wait for Clk_period;
		Addr <=  "0100110010010";
		Trees_din <= x"c1fee530";
		wait for Clk_period;
		Addr <=  "0100110010011";
		Trees_din <= x"83ffbd20";
		wait for Clk_period;
		Addr <=  "0100110010100";
		Trees_din <= x"1eff4a10";
		wait for Clk_period;
		Addr <=  "0100110010101";
		Trees_din <= x"baffeb08";
		wait for Clk_period;
		Addr <=  "0100110010110";
		Trees_din <= x"23ffa404";
		wait for Clk_period;
		Addr <=  "0100110010111";
		Trees_din <= x"ff7426fd";
		wait for Clk_period;
		Addr <=  "0100110011000";
		Trees_din <= x"001c26fd";
		wait for Clk_period;
		Addr <=  "0100110011001";
		Trees_din <= x"d3fed404";
		wait for Clk_period;
		Addr <=  "0100110011010";
		Trees_din <= x"ffdc26fd";
		wait for Clk_period;
		Addr <=  "0100110011011";
		Trees_din <= x"00ab26fd";
		wait for Clk_period;
		Addr <=  "0100110011100";
		Trees_din <= x"39000e08";
		wait for Clk_period;
		Addr <=  "0100110011101";
		Trees_din <= x"25ff7c04";
		wait for Clk_period;
		Addr <=  "0100110011110";
		Trees_din <= x"004126fd";
		wait for Clk_period;
		Addr <=  "0100110011111";
		Trees_din <= x"ff6e26fd";
		wait for Clk_period;
		Addr <=  "0100110100000";
		Trees_din <= x"09ffd204";
		wait for Clk_period;
		Addr <=  "0100110100001";
		Trees_din <= x"ff9526fd";
		wait for Clk_period;
		Addr <=  "0100110100010";
		Trees_din <= x"002a26fd";
		wait for Clk_period;
		Addr <=  "0100110100011";
		Trees_din <= x"7efeba08";
		wait for Clk_period;
		Addr <=  "0100110100100";
		Trees_din <= x"e5fefa04";
		wait for Clk_period;
		Addr <=  "0100110100101";
		Trees_din <= x"009a26fd";
		wait for Clk_period;
		Addr <=  "0100110100110";
		Trees_din <= x"fff326fd";
		wait for Clk_period;
		Addr <=  "0100110100111";
		Trees_din <= x"82ff4a04";
		wait for Clk_period;
		Addr <=  "0100110101000";
		Trees_din <= x"ff9826fd";
		wait for Clk_period;
		Addr <=  "0100110101001";
		Trees_din <= x"003f26fd";
		wait for Clk_period;
		Addr <=  "0100110101010";
		Trees_din <= x"67ff9318";
		wait for Clk_period;
		Addr <=  "0100110101011";
		Trees_din <= x"f1ff8608";
		wait for Clk_period;
		Addr <=  "0100110101100";
		Trees_din <= x"e3fea604";
		wait for Clk_period;
		Addr <=  "0100110101101";
		Trees_din <= x"fffa26fd";
		wait for Clk_period;
		Addr <=  "0100110101110";
		Trees_din <= x"ff6926fd";
		wait for Clk_period;
		Addr <=  "0100110101111";
		Trees_din <= x"c5ff3608";
		wait for Clk_period;
		Addr <=  "0100110110000";
		Trees_din <= x"d3feba04";
		wait for Clk_period;
		Addr <=  "0100110110001";
		Trees_din <= x"ffda26fd";
		wait for Clk_period;
		Addr <=  "0100110110010";
		Trees_din <= x"008626fd";
		wait for Clk_period;
		Addr <=  "0100110110011";
		Trees_din <= x"1b000d04";
		wait for Clk_period;
		Addr <=  "0100110110100";
		Trees_din <= x"ff9126fd";
		wait for Clk_period;
		Addr <=  "0100110110101";
		Trees_din <= x"002b26fd";
		wait for Clk_period;
		Addr <=  "0100110110110";
		Trees_din <= x"05003704";
		wait for Clk_period;
		Addr <=  "0100110110111";
		Trees_din <= x"ffb426fd";
		wait for Clk_period;
		Addr <=  "0100110111000";
		Trees_din <= x"7cfff108";
		wait for Clk_period;
		Addr <=  "0100110111001";
		Trees_din <= x"08006704";
		wait for Clk_period;
		Addr <=  "0100110111010";
		Trees_din <= x"002926fd";
		wait for Clk_period;
		Addr <=  "0100110111011";
		Trees_din <= x"00bc26fd";
		wait for Clk_period;
		Addr <=  "0100110111100";
		Trees_din <= x"b3ff2704";
		wait for Clk_period;
		Addr <=  "0100110111101";
		Trees_din <= x"006526fd";
		wait for Clk_period;
		Addr <=  "0100110111110";
		Trees_din <= x"ff9e26fd";
		wait for Clk_period;
		Addr <=  "0100110111111";
		Trees_din <= x"45ff1d4c";
		wait for Clk_period;
		Addr <=  "0100111000000";
		Trees_din <= x"d2ff9a3c";
		wait for Clk_period;
		Addr <=  "0100111000001";
		Trees_din <= x"00ffca20";
		wait for Clk_period;
		Addr <=  "0100111000010";
		Trees_din <= x"bcff8910";
		wait for Clk_period;
		Addr <=  "0100111000011";
		Trees_din <= x"3aff5708";
		wait for Clk_period;
		Addr <=  "0100111000100";
		Trees_din <= x"28ff2504";
		wait for Clk_period;
		Addr <=  "0100111000101";
		Trees_din <= x"001a2849";
		wait for Clk_period;
		Addr <=  "0100111000110";
		Trees_din <= x"ffea2849";
		wait for Clk_period;
		Addr <=  "0100111000111";
		Trees_din <= x"36fef404";
		wait for Clk_period;
		Addr <=  "0100111001000";
		Trees_din <= x"ffe52849";
		wait for Clk_period;
		Addr <=  "0100111001001";
		Trees_din <= x"00372849";
		wait for Clk_period;
		Addr <=  "0100111001010";
		Trees_din <= x"e1ffaa08";
		wait for Clk_period;
		Addr <=  "0100111001011";
		Trees_din <= x"09006704";
		wait for Clk_period;
		Addr <=  "0100111001100";
		Trees_din <= x"ff8d2849";
		wait for Clk_period;
		Addr <=  "0100111001101";
		Trees_din <= x"004c2849";
		wait for Clk_period;
		Addr <=  "0100111001110";
		Trees_din <= x"26003a04";
		wait for Clk_period;
		Addr <=  "0100111001111";
		Trees_din <= x"ffbb2849";
		wait for Clk_period;
		Addr <=  "0100111010000";
		Trees_din <= x"003b2849";
		wait for Clk_period;
		Addr <=  "0100111010001";
		Trees_din <= x"8cffaf0c";
		wait for Clk_period;
		Addr <=  "0100111010010";
		Trees_din <= x"c3ff4a04";
		wait for Clk_period;
		Addr <=  "0100111010011";
		Trees_din <= x"002d2849";
		wait for Clk_period;
		Addr <=  "0100111010100";
		Trees_din <= x"76005b04";
		wait for Clk_period;
		Addr <=  "0100111010101";
		Trees_din <= x"ff632849";
		wait for Clk_period;
		Addr <=  "0100111010110";
		Trees_din <= x"00072849";
		wait for Clk_period;
		Addr <=  "0100111010111";
		Trees_din <= x"f3fe9808";
		wait for Clk_period;
		Addr <=  "0100111011000";
		Trees_din <= x"2f000204";
		wait for Clk_period;
		Addr <=  "0100111011001";
		Trees_din <= x"007f2849";
		wait for Clk_period;
		Addr <=  "0100111011010";
		Trees_din <= x"ffdc2849";
		wait for Clk_period;
		Addr <=  "0100111011011";
		Trees_din <= x"a9ff3504";
		wait for Clk_period;
		Addr <=  "0100111011100";
		Trees_din <= x"00442849";
		wait for Clk_period;
		Addr <=  "0100111011101";
		Trees_din <= x"ffab2849";
		wait for Clk_period;
		Addr <=  "0100111011110";
		Trees_din <= x"30001d0c";
		wait for Clk_period;
		Addr <=  "0100111011111";
		Trees_din <= x"d8001e04";
		wait for Clk_period;
		Addr <=  "0100111100000";
		Trees_din <= x"ffef2849";
		wait for Clk_period;
		Addr <=  "0100111100001";
		Trees_din <= x"c3ffb604";
		wait for Clk_period;
		Addr <=  "0100111100010";
		Trees_din <= x"00352849";
		wait for Clk_period;
		Addr <=  "0100111100011";
		Trees_din <= x"00c62849";
		wait for Clk_period;
		Addr <=  "0100111100100";
		Trees_din <= x"ffc22849";
		wait for Clk_period;
		Addr <=  "0100111100101";
		Trees_din <= x"a5ff7138";
		wait for Clk_period;
		Addr <=  "0100111100110";
		Trees_din <= x"0800e920";
		wait for Clk_period;
		Addr <=  "0100111100111";
		Trees_din <= x"f1ff7210";
		wait for Clk_period;
		Addr <=  "0100111101000";
		Trees_din <= x"49ffe308";
		wait for Clk_period;
		Addr <=  "0100111101001";
		Trees_din <= x"5fff7a04";
		wait for Clk_period;
		Addr <=  "0100111101010";
		Trees_din <= x"00682849";
		wait for Clk_period;
		Addr <=  "0100111101011";
		Trees_din <= x"ffd02849";
		wait for Clk_period;
		Addr <=  "0100111101100";
		Trees_din <= x"b5fe5204";
		wait for Clk_period;
		Addr <=  "0100111101101";
		Trees_din <= x"00602849";
		wait for Clk_period;
		Addr <=  "0100111101110";
		Trees_din <= x"ffb02849";
		wait for Clk_period;
		Addr <=  "0100111101111";
		Trees_din <= x"bcfefd08";
		wait for Clk_period;
		Addr <=  "0100111110000";
		Trees_din <= x"77feaa04";
		wait for Clk_period;
		Addr <=  "0100111110001";
		Trees_din <= x"00542849";
		wait for Clk_period;
		Addr <=  "0100111110010";
		Trees_din <= x"ffd62849";
		wait for Clk_period;
		Addr <=  "0100111110011";
		Trees_din <= x"71001b04";
		wait for Clk_period;
		Addr <=  "0100111110100";
		Trees_din <= x"ffaa2849";
		wait for Clk_period;
		Addr <=  "0100111110101";
		Trees_din <= x"00492849";
		wait for Clk_period;
		Addr <=  "0100111110110";
		Trees_din <= x"5cffce08";
		wait for Clk_period;
		Addr <=  "0100111110111";
		Trees_din <= x"27ffb604";
		wait for Clk_period;
		Addr <=  "0100111111000";
		Trees_din <= x"fff42849";
		wait for Clk_period;
		Addr <=  "0100111111001";
		Trees_din <= x"ff892849";
		wait for Clk_period;
		Addr <=  "0100111111010";
		Trees_din <= x"73ffb908";
		wait for Clk_period;
		Addr <=  "0100111111011";
		Trees_din <= x"2bffab04";
		wait for Clk_period;
		Addr <=  "0100111111100";
		Trees_din <= x"00362849";
		wait for Clk_period;
		Addr <=  "0100111111101";
		Trees_din <= x"ff8e2849";
		wait for Clk_period;
		Addr <=  "0100111111110";
		Trees_din <= x"1fffcc04";
		wait for Clk_period;
		Addr <=  "0100111111111";
		Trees_din <= x"ffef2849";
		wait for Clk_period;
		Addr <=  "0101000000000";
		Trees_din <= x"00972849";
		wait for Clk_period;
		Addr <=  "0101000000001";
		Trees_din <= x"e4fe8810";
		wait for Clk_period;
		Addr <=  "0101000000010";
		Trees_din <= x"67ffb008";
		wait for Clk_period;
		Addr <=  "0101000000011";
		Trees_din <= x"8cff4004";
		wait for Clk_period;
		Addr <=  "0101000000100";
		Trees_din <= x"00162849";
		wait for Clk_period;
		Addr <=  "0101000000101";
		Trees_din <= x"ff732849";
		wait for Clk_period;
		Addr <=  "0101000000110";
		Trees_din <= x"de005604";
		wait for Clk_period;
		Addr <=  "0101000000111";
		Trees_din <= x"fff62849";
		wait for Clk_period;
		Addr <=  "0101000001000";
		Trees_din <= x"007c2849";
		wait for Clk_period;
		Addr <=  "0101000001001";
		Trees_din <= x"59ff0808";
		wait for Clk_period;
		Addr <=  "0101000001010";
		Trees_din <= x"a8ff5804";
		wait for Clk_period;
		Addr <=  "0101000001011";
		Trees_din <= x"00332849";
		wait for Clk_period;
		Addr <=  "0101000001100";
		Trees_din <= x"ff8a2849";
		wait for Clk_period;
		Addr <=  "0101000001101";
		Trees_din <= x"99fe8504";
		wait for Clk_period;
		Addr <=  "0101000001110";
		Trees_din <= x"ffbd2849";
		wait for Clk_period;
		Addr <=  "0101000001111";
		Trees_din <= x"72fffa04";
		wait for Clk_period;
		Addr <=  "0101000010000";
		Trees_din <= x"00312849";
		wait for Clk_period;
		Addr <=  "0101000010001";
		Trees_din <= x"00a52849";
		wait for Clk_period;
		Addr <=  "0101000010010";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0101000010011";
		Trees_din <= x"dcfe6518";
		wait for Clk_period;
		Addr <=  "0101000010100";
		Trees_din <= x"65ffbd14";
		wait for Clk_period;
		Addr <=  "0101000010101";
		Trees_din <= x"6d003e0c";
		wait for Clk_period;
		Addr <=  "0101000010110";
		Trees_din <= x"65ff3f04";
		wait for Clk_period;
		Addr <=  "0101000010111";
		Trees_din <= x"00842951";
		wait for Clk_period;
		Addr <=  "0101000011000";
		Trees_din <= x"d3ff1704";
		wait for Clk_period;
		Addr <=  "0101000011001";
		Trees_din <= x"ff882951";
		wait for Clk_period;
		Addr <=  "0101000011010";
		Trees_din <= x"00142951";
		wait for Clk_period;
		Addr <=  "0101000011011";
		Trees_din <= x"5bff4704";
		wait for Clk_period;
		Addr <=  "0101000011100";
		Trees_din <= x"00202951";
		wait for Clk_period;
		Addr <=  "0101000011101";
		Trees_din <= x"00b42951";
		wait for Clk_period;
		Addr <=  "0101000011110";
		Trees_din <= x"ff962951";
		wait for Clk_period;
		Addr <=  "0101000011111";
		Trees_din <= x"cdffe540";
		wait for Clk_period;
		Addr <=  "0101000100000";
		Trees_din <= x"adffae20";
		wait for Clk_period;
		Addr <=  "0101000100001";
		Trees_din <= x"40ffb910";
		wait for Clk_period;
		Addr <=  "0101000100010";
		Trees_din <= x"0eff6408";
		wait for Clk_period;
		Addr <=  "0101000100011";
		Trees_din <= x"95feb704";
		wait for Clk_period;
		Addr <=  "0101000100100";
		Trees_din <= x"003c2951";
		wait for Clk_period;
		Addr <=  "0101000100101";
		Trees_din <= x"ff852951";
		wait for Clk_period;
		Addr <=  "0101000100110";
		Trees_din <= x"b2001304";
		wait for Clk_period;
		Addr <=  "0101000100111";
		Trees_din <= x"000f2951";
		wait for Clk_period;
		Addr <=  "0101000101000";
		Trees_din <= x"00902951";
		wait for Clk_period;
		Addr <=  "0101000101001";
		Trees_din <= x"de008f08";
		wait for Clk_period;
		Addr <=  "0101000101010";
		Trees_din <= x"efff5604";
		wait for Clk_period;
		Addr <=  "0101000101011";
		Trees_din <= x"ffdb2951";
		wait for Clk_period;
		Addr <=  "0101000101100";
		Trees_din <= x"00102951";
		wait for Clk_period;
		Addr <=  "0101000101101";
		Trees_din <= x"84000204";
		wait for Clk_period;
		Addr <=  "0101000101110";
		Trees_din <= x"00522951";
		wait for Clk_period;
		Addr <=  "0101000101111";
		Trees_din <= x"ffb12951";
		wait for Clk_period;
		Addr <=  "0101000110000";
		Trees_din <= x"45fe6010";
		wait for Clk_period;
		Addr <=  "0101000110001";
		Trees_din <= x"eeff9008";
		wait for Clk_period;
		Addr <=  "0101000110010";
		Trees_din <= x"b0ff4a04";
		wait for Clk_period;
		Addr <=  "0101000110011";
		Trees_din <= x"ffd92951";
		wait for Clk_period;
		Addr <=  "0101000110100";
		Trees_din <= x"006f2951";
		wait for Clk_period;
		Addr <=  "0101000110101";
		Trees_din <= x"77ff5904";
		wait for Clk_period;
		Addr <=  "0101000110110";
		Trees_din <= x"ff6f2951";
		wait for Clk_period;
		Addr <=  "0101000110111";
		Trees_din <= x"000f2951";
		wait for Clk_period;
		Addr <=  "0101000111000";
		Trees_din <= x"68fe1008";
		wait for Clk_period;
		Addr <=  "0101000111001";
		Trees_din <= x"ab002604";
		wait for Clk_period;
		Addr <=  "0101000111010";
		Trees_din <= x"fff32951";
		wait for Clk_period;
		Addr <=  "0101000111011";
		Trees_din <= x"ff7c2951";
		wait for Clk_period;
		Addr <=  "0101000111100";
		Trees_din <= x"43ff4f04";
		wait for Clk_period;
		Addr <=  "0101000111101";
		Trees_din <= x"00562951";
		wait for Clk_period;
		Addr <=  "0101000111110";
		Trees_din <= x"00192951";
		wait for Clk_period;
		Addr <=  "0101000111111";
		Trees_din <= x"8c010c20";
		wait for Clk_period;
		Addr <=  "0101001000000";
		Trees_din <= x"f3fe5a10";
		wait for Clk_period;
		Addr <=  "0101001000001";
		Trees_din <= x"39ff8908";
		wait for Clk_period;
		Addr <=  "0101001000010";
		Trees_din <= x"12ffa904";
		wait for Clk_period;
		Addr <=  "0101001000011";
		Trees_din <= x"ff732951";
		wait for Clk_period;
		Addr <=  "0101001000100";
		Trees_din <= x"00152951";
		wait for Clk_period;
		Addr <=  "0101001000101";
		Trees_din <= x"d3fec104";
		wait for Clk_period;
		Addr <=  "0101001000110";
		Trees_din <= x"ffba2951";
		wait for Clk_period;
		Addr <=  "0101001000111";
		Trees_din <= x"006e2951";
		wait for Clk_period;
		Addr <=  "0101001001000";
		Trees_din <= x"05005e08";
		wait for Clk_period;
		Addr <=  "0101001001001";
		Trees_din <= x"edff4504";
		wait for Clk_period;
		Addr <=  "0101001001010";
		Trees_din <= x"00372951";
		wait for Clk_period;
		Addr <=  "0101001001011";
		Trees_din <= x"ffc12951";
		wait for Clk_period;
		Addr <=  "0101001001100";
		Trees_din <= x"dfff1504";
		wait for Clk_period;
		Addr <=  "0101001001101";
		Trees_din <= x"ffb42951";
		wait for Clk_period;
		Addr <=  "0101001001110";
		Trees_din <= x"000f2951";
		wait for Clk_period;
		Addr <=  "0101001001111";
		Trees_din <= x"db00a404";
		wait for Clk_period;
		Addr <=  "0101001010000";
		Trees_din <= x"008a2951";
		wait for Clk_period;
		Addr <=  "0101001010001";
		Trees_din <= x"9affa204";
		wait for Clk_period;
		Addr <=  "0101001010010";
		Trees_din <= x"ffab2951";
		wait for Clk_period;
		Addr <=  "0101001010011";
		Trees_din <= x"00422951";
		wait for Clk_period;
		Addr <=  "0101001010100";
		Trees_din <= x"7efdfc28";
		wait for Clk_period;
		Addr <=  "0101001010101";
		Trees_din <= x"daff1804";
		wait for Clk_period;
		Addr <=  "0101001010110";
		Trees_din <= x"ff8d2a8d";
		wait for Clk_period;
		Addr <=  "0101001010111";
		Trees_din <= x"2e000a18";
		wait for Clk_period;
		Addr <=  "0101001011000";
		Trees_din <= x"67fed10c";
		wait for Clk_period;
		Addr <=  "0101001011001";
		Trees_din <= x"5c005e04";
		wait for Clk_period;
		Addr <=  "0101001011010";
		Trees_din <= x"ff9b2a8d";
		wait for Clk_period;
		Addr <=  "0101001011011";
		Trees_din <= x"adff8104";
		wait for Clk_period;
		Addr <=  "0101001011100";
		Trees_din <= x"ffe22a8d";
		wait for Clk_period;
		Addr <=  "0101001011101";
		Trees_din <= x"00622a8d";
		wait for Clk_period;
		Addr <=  "0101001011110";
		Trees_din <= x"7afede04";
		wait for Clk_period;
		Addr <=  "0101001011111";
		Trees_din <= x"ffb42a8d";
		wait for Clk_period;
		Addr <=  "0101001100000";
		Trees_din <= x"3bfedf04";
		wait for Clk_period;
		Addr <=  "0101001100001";
		Trees_din <= x"ffd42a8d";
		wait for Clk_period;
		Addr <=  "0101001100010";
		Trees_din <= x"00842a8d";
		wait for Clk_period;
		Addr <=  "0101001100011";
		Trees_din <= x"ac006b08";
		wait for Clk_period;
		Addr <=  "0101001100100";
		Trees_din <= x"69ff4104";
		wait for Clk_period;
		Addr <=  "0101001100101";
		Trees_din <= x"ffeb2a8d";
		wait for Clk_period;
		Addr <=  "0101001100110";
		Trees_din <= x"ff852a8d";
		wait for Clk_period;
		Addr <=  "0101001100111";
		Trees_din <= x"003f2a8d";
		wait for Clk_period;
		Addr <=  "0101001101000";
		Trees_din <= x"b1ff4c3c";
		wait for Clk_period;
		Addr <=  "0101001101001";
		Trees_din <= x"7400011c";
		wait for Clk_period;
		Addr <=  "0101001101010";
		Trees_din <= x"8fff6910";
		wait for Clk_period;
		Addr <=  "0101001101011";
		Trees_din <= x"81ff3908";
		wait for Clk_period;
		Addr <=  "0101001101100";
		Trees_din <= x"c3fff104";
		wait for Clk_period;
		Addr <=  "0101001101101";
		Trees_din <= x"fff12a8d";
		wait for Clk_period;
		Addr <=  "0101001101110";
		Trees_din <= x"005d2a8d";
		wait for Clk_period;
		Addr <=  "0101001101111";
		Trees_din <= x"36ffc904";
		wait for Clk_period;
		Addr <=  "0101001110000";
		Trees_din <= x"ffef2a8d";
		wait for Clk_period;
		Addr <=  "0101001110001";
		Trees_din <= x"00332a8d";
		wait for Clk_period;
		Addr <=  "0101001110010";
		Trees_din <= x"b1ff4308";
		wait for Clk_period;
		Addr <=  "0101001110011";
		Trees_din <= x"46fed304";
		wait for Clk_period;
		Addr <=  "0101001110100";
		Trees_din <= x"fff02a8d";
		wait for Clk_period;
		Addr <=  "0101001110101";
		Trees_din <= x"006f2a8d";
		wait for Clk_period;
		Addr <=  "0101001110110";
		Trees_din <= x"ff862a8d";
		wait for Clk_period;
		Addr <=  "0101001110111";
		Trees_din <= x"99fe5510";
		wait for Clk_period;
		Addr <=  "0101001111000";
		Trees_din <= x"92ff4508";
		wait for Clk_period;
		Addr <=  "0101001111001";
		Trees_din <= x"0aff8004";
		wait for Clk_period;
		Addr <=  "0101001111010";
		Trees_din <= x"ff882a8d";
		wait for Clk_period;
		Addr <=  "0101001111011";
		Trees_din <= x"005a2a8d";
		wait for Clk_period;
		Addr <=  "0101001111100";
		Trees_din <= x"56fff104";
		wait for Clk_period;
		Addr <=  "0101001111101";
		Trees_din <= x"ff802a8d";
		wait for Clk_period;
		Addr <=  "0101001111110";
		Trees_din <= x"00702a8d";
		wait for Clk_period;
		Addr <=  "0101001111111";
		Trees_din <= x"40006308";
		wait for Clk_period;
		Addr <=  "0101010000000";
		Trees_din <= x"3dff4a04";
		wait for Clk_period;
		Addr <=  "0101010000001";
		Trees_din <= x"004a2a8d";
		wait for Clk_period;
		Addr <=  "0101010000010";
		Trees_din <= x"ffc32a8d";
		wait for Clk_period;
		Addr <=  "0101010000011";
		Trees_din <= x"ab006404";
		wait for Clk_period;
		Addr <=  "0101010000100";
		Trees_din <= x"00502a8d";
		wait for Clk_period;
		Addr <=  "0101010000101";
		Trees_din <= x"ffca2a8d";
		wait for Clk_period;
		Addr <=  "0101010000110";
		Trees_din <= x"f1ff931c";
		wait for Clk_period;
		Addr <=  "0101010000111";
		Trees_din <= x"b9fe5b0c";
		wait for Clk_period;
		Addr <=  "0101010001000";
		Trees_din <= x"3ffff104";
		wait for Clk_period;
		Addr <=  "0101010001001";
		Trees_din <= x"ff792a8d";
		wait for Clk_period;
		Addr <=  "0101010001010";
		Trees_din <= x"45fedf04";
		wait for Clk_period;
		Addr <=  "0101010001011";
		Trees_din <= x"00502a8d";
		wait for Clk_period;
		Addr <=  "0101010001100";
		Trees_din <= x"ffa62a8d";
		wait for Clk_period;
		Addr <=  "0101010001101";
		Trees_din <= x"a1ffcc08";
		wait for Clk_period;
		Addr <=  "0101010001110";
		Trees_din <= x"70fe3304";
		wait for Clk_period;
		Addr <=  "0101010001111";
		Trees_din <= x"ff962a8d";
		wait for Clk_period;
		Addr <=  "0101010010000";
		Trees_din <= x"00562a8d";
		wait for Clk_period;
		Addr <=  "0101010010001";
		Trees_din <= x"d0003204";
		wait for Clk_period;
		Addr <=  "0101010010010";
		Trees_din <= x"00482a8d";
		wait for Clk_period;
		Addr <=  "0101010010011";
		Trees_din <= x"ff922a8d";
		wait for Clk_period;
		Addr <=  "0101010010100";
		Trees_din <= x"b3ff7810";
		wait for Clk_period;
		Addr <=  "0101010010101";
		Trees_din <= x"6d003d08";
		wait for Clk_period;
		Addr <=  "0101010010110";
		Trees_din <= x"9dff9404";
		wait for Clk_period;
		Addr <=  "0101010010111";
		Trees_din <= x"fff12a8d";
		wait for Clk_period;
		Addr <=  "0101010011000";
		Trees_din <= x"ff812a8d";
		wait for Clk_period;
		Addr <=  "0101010011001";
		Trees_din <= x"bfff4d04";
		wait for Clk_period;
		Addr <=  "0101010011010";
		Trees_din <= x"004b2a8d";
		wait for Clk_period;
		Addr <=  "0101010011011";
		Trees_din <= x"ffdc2a8d";
		wait for Clk_period;
		Addr <=  "0101010011100";
		Trees_din <= x"5dffe908";
		wait for Clk_period;
		Addr <=  "0101010011101";
		Trees_din <= x"1effea04";
		wait for Clk_period;
		Addr <=  "0101010011110";
		Trees_din <= x"00a42a8d";
		wait for Clk_period;
		Addr <=  "0101010011111";
		Trees_din <= x"ffea2a8d";
		wait for Clk_period;
		Addr <=  "0101010100000";
		Trees_din <= x"99fe9004";
		wait for Clk_period;
		Addr <=  "0101010100001";
		Trees_din <= x"00762a8d";
		wait for Clk_period;
		Addr <=  "0101010100010";
		Trees_din <= x"ffa92a8d";
		wait for Clk_period;
		Addr <=  "0101010100011";
		Trees_din <= x"2eff3558";
		wait for Clk_period;
		Addr <=  "0101010100100";
		Trees_din <= x"6fffcb38";
		wait for Clk_period;
		Addr <=  "0101010100101";
		Trees_din <= x"9bff6820";
		wait for Clk_period;
		Addr <=  "0101010100110";
		Trees_din <= x"65ff8710";
		wait for Clk_period;
		Addr <=  "0101010100111";
		Trees_din <= x"c7ff7e08";
		wait for Clk_period;
		Addr <=  "0101010101000";
		Trees_din <= x"89008204";
		wait for Clk_period;
		Addr <=  "0101010101001";
		Trees_din <= x"007a2c21";
		wait for Clk_period;
		Addr <=  "0101010101010";
		Trees_din <= x"ffde2c21";
		wait for Clk_period;
		Addr <=  "0101010101011";
		Trees_din <= x"e5fedb04";
		wait for Clk_period;
		Addr <=  "0101010101100";
		Trees_din <= x"ff8e2c21";
		wait for Clk_period;
		Addr <=  "0101010101101";
		Trees_din <= x"001a2c21";
		wait for Clk_period;
		Addr <=  "0101010101110";
		Trees_din <= x"c9ffad08";
		wait for Clk_period;
		Addr <=  "0101010101111";
		Trees_din <= x"60ff8204";
		wait for Clk_period;
		Addr <=  "0101010110000";
		Trees_din <= x"ffa12c21";
		wait for Clk_period;
		Addr <=  "0101010110001";
		Trees_din <= x"007c2c21";
		wait for Clk_period;
		Addr <=  "0101010110010";
		Trees_din <= x"93ffdf04";
		wait for Clk_period;
		Addr <=  "0101010110011";
		Trees_din <= x"ff752c21";
		wait for Clk_period;
		Addr <=  "0101010110100";
		Trees_din <= x"001e2c21";
		wait for Clk_period;
		Addr <=  "0101010110101";
		Trees_din <= x"a6000610";
		wait for Clk_period;
		Addr <=  "0101010110110";
		Trees_din <= x"eaff6a08";
		wait for Clk_period;
		Addr <=  "0101010110111";
		Trees_din <= x"81ffe004";
		wait for Clk_period;
		Addr <=  "0101010111000";
		Trees_din <= x"ffb42c21";
		wait for Clk_period;
		Addr <=  "0101010111001";
		Trees_din <= x"00472c21";
		wait for Clk_period;
		Addr <=  "0101010111010";
		Trees_din <= x"39003904";
		wait for Clk_period;
		Addr <=  "0101010111011";
		Trees_din <= x"ff712c21";
		wait for Clk_period;
		Addr <=  "0101010111100";
		Trees_din <= x"ffe62c21";
		wait for Clk_period;
		Addr <=  "0101010111101";
		Trees_din <= x"4eff9b04";
		wait for Clk_period;
		Addr <=  "0101010111110";
		Trees_din <= x"000d2c21";
		wait for Clk_period;
		Addr <=  "0101010111111";
		Trees_din <= x"00792c21";
		wait for Clk_period;
		Addr <=  "0101011000000";
		Trees_din <= x"daffcc0c";
		wait for Clk_period;
		Addr <=  "0101011000001";
		Trees_din <= x"30ff7204";
		wait for Clk_period;
		Addr <=  "0101011000010";
		Trees_din <= x"006c2c21";
		wait for Clk_period;
		Addr <=  "0101011000011";
		Trees_din <= x"d1ff1a04";
		wait for Clk_period;
		Addr <=  "0101011000100";
		Trees_din <= x"002d2c21";
		wait for Clk_period;
		Addr <=  "0101011000101";
		Trees_din <= x"ff832c21";
		wait for Clk_period;
		Addr <=  "0101011000110";
		Trees_din <= x"cafdbf08";
		wait for Clk_period;
		Addr <=  "0101011000111";
		Trees_din <= x"f0ffb704";
		wait for Clk_period;
		Addr <=  "0101011001000";
		Trees_din <= x"ffb22c21";
		wait for Clk_period;
		Addr <=  "0101011001001";
		Trees_din <= x"00582c21";
		wait for Clk_period;
		Addr <=  "0101011001010";
		Trees_din <= x"d4ffd808";
		wait for Clk_period;
		Addr <=  "0101011001011";
		Trees_din <= x"21ffec04";
		wait for Clk_period;
		Addr <=  "0101011001100";
		Trees_din <= x"00a92c21";
		wait for Clk_period;
		Addr <=  "0101011001101";
		Trees_din <= x"00242c21";
		wait for Clk_period;
		Addr <=  "0101011001110";
		Trees_din <= x"fff42c21";
		wait for Clk_period;
		Addr <=  "0101011001111";
		Trees_din <= x"aeff433c";
		wait for Clk_period;
		Addr <=  "0101011010000";
		Trees_din <= x"55008320";
		wait for Clk_period;
		Addr <=  "0101011010001";
		Trees_din <= x"b1ff3510";
		wait for Clk_period;
		Addr <=  "0101011010010";
		Trees_din <= x"98ff1408";
		wait for Clk_period;
		Addr <=  "0101011010011";
		Trees_din <= x"68ff3c04";
		wait for Clk_period;
		Addr <=  "0101011010100";
		Trees_din <= x"001a2c21";
		wait for Clk_period;
		Addr <=  "0101011010101";
		Trees_din <= x"ffd42c21";
		wait for Clk_period;
		Addr <=  "0101011010110";
		Trees_din <= x"ec004404";
		wait for Clk_period;
		Addr <=  "0101011010111";
		Trees_din <= x"ffd62c21";
		wait for Clk_period;
		Addr <=  "0101011011000";
		Trees_din <= x"00382c21";
		wait for Clk_period;
		Addr <=  "0101011011001";
		Trees_din <= x"3bff5008";
		wait for Clk_period;
		Addr <=  "0101011011010";
		Trees_din <= x"67fff104";
		wait for Clk_period;
		Addr <=  "0101011011011";
		Trees_din <= x"000f2c21";
		wait for Clk_period;
		Addr <=  "0101011011100";
		Trees_din <= x"ff7b2c21";
		wait for Clk_period;
		Addr <=  "0101011011101";
		Trees_din <= x"62ff3604";
		wait for Clk_period;
		Addr <=  "0101011011110";
		Trees_din <= x"00702c21";
		wait for Clk_period;
		Addr <=  "0101011011111";
		Trees_din <= x"001a2c21";
		wait for Clk_period;
		Addr <=  "0101011100000";
		Trees_din <= x"bbff560c";
		wait for Clk_period;
		Addr <=  "0101011100001";
		Trees_din <= x"72009308";
		wait for Clk_period;
		Addr <=  "0101011100010";
		Trees_din <= x"3bfefe04";
		wait for Clk_period;
		Addr <=  "0101011100011";
		Trees_din <= x"000a2c21";
		wait for Clk_period;
		Addr <=  "0101011100100";
		Trees_din <= x"ff8c2c21";
		wait for Clk_period;
		Addr <=  "0101011100101";
		Trees_din <= x"00552c21";
		wait for Clk_period;
		Addr <=  "0101011100110";
		Trees_din <= x"c1fee308";
		wait for Clk_period;
		Addr <=  "0101011100111";
		Trees_din <= x"efff2504";
		wait for Clk_period;
		Addr <=  "0101011101000";
		Trees_din <= x"00712c21";
		wait for Clk_period;
		Addr <=  "0101011101001";
		Trees_din <= x"ffb42c21";
		wait for Clk_period;
		Addr <=  "0101011101010";
		Trees_din <= x"17ffdb04";
		wait for Clk_period;
		Addr <=  "0101011101011";
		Trees_din <= x"ffe02c21";
		wait for Clk_period;
		Addr <=  "0101011101100";
		Trees_din <= x"008a2c21";
		wait for Clk_period;
		Addr <=  "0101011101101";
		Trees_din <= x"9bfed618";
		wait for Clk_period;
		Addr <=  "0101011101110";
		Trees_din <= x"a1fec308";
		wait for Clk_period;
		Addr <=  "0101011101111";
		Trees_din <= x"3f000704";
		wait for Clk_period;
		Addr <=  "0101011110000";
		Trees_din <= x"ff7f2c21";
		wait for Clk_period;
		Addr <=  "0101011110001";
		Trees_din <= x"fffa2c21";
		wait for Clk_period;
		Addr <=  "0101011110010";
		Trees_din <= x"22ffd708";
		wait for Clk_period;
		Addr <=  "0101011110011";
		Trees_din <= x"b8ff1e04";
		wait for Clk_period;
		Addr <=  "0101011110100";
		Trees_din <= x"00392c21";
		wait for Clk_period;
		Addr <=  "0101011110101";
		Trees_din <= x"ff912c21";
		wait for Clk_period;
		Addr <=  "0101011110110";
		Trees_din <= x"d5ffc404";
		wait for Clk_period;
		Addr <=  "0101011110111";
		Trees_din <= x"ffd52c21";
		wait for Clk_period;
		Addr <=  "0101011111000";
		Trees_din <= x"00872c21";
		wait for Clk_period;
		Addr <=  "0101011111001";
		Trees_din <= x"86ff1a10";
		wait for Clk_period;
		Addr <=  "0101011111010";
		Trees_din <= x"41ff4008";
		wait for Clk_period;
		Addr <=  "0101011111011";
		Trees_din <= x"b6ff8504";
		wait for Clk_period;
		Addr <=  "0101011111100";
		Trees_din <= x"ffee2c21";
		wait for Clk_period;
		Addr <=  "0101011111101";
		Trees_din <= x"00502c21";
		wait for Clk_period;
		Addr <=  "0101011111110";
		Trees_din <= x"5fffdc04";
		wait for Clk_period;
		Addr <=  "0101011111111";
		Trees_din <= x"ff8e2c21";
		wait for Clk_period;
		Addr <=  "0101100000000";
		Trees_din <= x"00622c21";
		wait for Clk_period;
		Addr <=  "0101100000001";
		Trees_din <= x"f5ffb908";
		wait for Clk_period;
		Addr <=  "0101100000010";
		Trees_din <= x"dcff7004";
		wait for Clk_period;
		Addr <=  "0101100000011";
		Trees_din <= x"00842c21";
		wait for Clk_period;
		Addr <=  "0101100000100";
		Trees_din <= x"ffc52c21";
		wait for Clk_period;
		Addr <=  "0101100000101";
		Trees_din <= x"e2ffb804";
		wait for Clk_period;
		Addr <=  "0101100000110";
		Trees_din <= x"ff832c21";
		wait for Clk_period;
		Addr <=  "0101100000111";
		Trees_din <= x"00022c21";
		wait for Clk_period;
		Addr <=  "0101100001000";
		Trees_din <= x"44005368";
		wait for Clk_period;
		Addr <=  "0101100001001";
		Trees_din <= x"0700b134";
		wait for Clk_period;
		Addr <=  "0101100001010";
		Trees_din <= x"c800a220";
		wait for Clk_period;
		Addr <=  "0101100001011";
		Trees_din <= x"83ff1510";
		wait for Clk_period;
		Addr <=  "0101100001100";
		Trees_din <= x"33feea08";
		wait for Clk_period;
		Addr <=  "0101100001101";
		Trees_din <= x"70fe8604";
		wait for Clk_period;
		Addr <=  "0101100001110";
		Trees_din <= x"ffc82d65";
		wait for Clk_period;
		Addr <=  "0101100001111";
		Trees_din <= x"002f2d65";
		wait for Clk_period;
		Addr <=  "0101100010000";
		Trees_din <= x"8e00cb04";
		wait for Clk_period;
		Addr <=  "0101100010001";
		Trees_din <= x"ffba2d65";
		wait for Clk_period;
		Addr <=  "0101100010010";
		Trees_din <= x"00562d65";
		wait for Clk_period;
		Addr <=  "0101100010011";
		Trees_din <= x"d1ff5808";
		wait for Clk_period;
		Addr <=  "0101100010100";
		Trees_din <= x"15ff4704";
		wait for Clk_period;
		Addr <=  "0101100010101";
		Trees_din <= x"ffc52d65";
		wait for Clk_period;
		Addr <=  "0101100010110";
		Trees_din <= x"00022d65";
		wait for Clk_period;
		Addr <=  "0101100010111";
		Trees_din <= x"c4ffc904";
		wait for Clk_period;
		Addr <=  "0101100011000";
		Trees_din <= x"00112d65";
		wait for Clk_period;
		Addr <=  "0101100011001";
		Trees_din <= x"008a2d65";
		wait for Clk_period;
		Addr <=  "0101100011010";
		Trees_din <= x"ccff6f08";
		wait for Clk_period;
		Addr <=  "0101100011011";
		Trees_din <= x"22000104";
		wait for Clk_period;
		Addr <=  "0101100011100";
		Trees_din <= x"00102d65";
		wait for Clk_period;
		Addr <=  "0101100011101";
		Trees_din <= x"ff8c2d65";
		wait for Clk_period;
		Addr <=  "0101100011110";
		Trees_din <= x"9a004f08";
		wait for Clk_period;
		Addr <=  "0101100011111";
		Trees_din <= x"58ff1504";
		wait for Clk_period;
		Addr <=  "0101100100000";
		Trees_din <= x"009b2d65";
		wait for Clk_period;
		Addr <=  "0101100100001";
		Trees_din <= x"ffed2d65";
		wait for Clk_period;
		Addr <=  "0101100100010";
		Trees_din <= x"ffbb2d65";
		wait for Clk_period;
		Addr <=  "0101100100011";
		Trees_din <= x"e6fff820";
		wait for Clk_period;
		Addr <=  "0101100100100";
		Trees_din <= x"f9ff6e10";
		wait for Clk_period;
		Addr <=  "0101100100101";
		Trees_din <= x"7dffb008";
		wait for Clk_period;
		Addr <=  "0101100100110";
		Trees_din <= x"8b006004";
		wait for Clk_period;
		Addr <=  "0101100100111";
		Trees_din <= x"00522d65";
		wait for Clk_period;
		Addr <=  "0101100101000";
		Trees_din <= x"ffa02d65";
		wait for Clk_period;
		Addr <=  "0101100101001";
		Trees_din <= x"53ff9504";
		wait for Clk_period;
		Addr <=  "0101100101010";
		Trees_din <= x"ffdc2d65";
		wait for Clk_period;
		Addr <=  "0101100101011";
		Trees_din <= x"00292d65";
		wait for Clk_period;
		Addr <=  "0101100101100";
		Trees_din <= x"d9ff8108";
		wait for Clk_period;
		Addr <=  "0101100101101";
		Trees_din <= x"3d002404";
		wait for Clk_period;
		Addr <=  "0101100101110";
		Trees_din <= x"006e2d65";
		wait for Clk_period;
		Addr <=  "0101100101111";
		Trees_din <= x"ffcc2d65";
		wait for Clk_period;
		Addr <=  "0101100110000";
		Trees_din <= x"1efefb04";
		wait for Clk_period;
		Addr <=  "0101100110001";
		Trees_din <= x"00432d65";
		wait for Clk_period;
		Addr <=  "0101100110010";
		Trees_din <= x"ff9f2d65";
		wait for Clk_period;
		Addr <=  "0101100110011";
		Trees_din <= x"94feec08";
		wait for Clk_period;
		Addr <=  "0101100110100";
		Trees_din <= x"efff7f04";
		wait for Clk_period;
		Addr <=  "0101100110101";
		Trees_din <= x"00082d65";
		wait for Clk_period;
		Addr <=  "0101100110110";
		Trees_din <= x"ffa32d65";
		wait for Clk_period;
		Addr <=  "0101100110111";
		Trees_din <= x"37ffe708";
		wait for Clk_period;
		Addr <=  "0101100111000";
		Trees_din <= x"00ffaa04";
		wait for Clk_period;
		Addr <=  "0101100111001";
		Trees_din <= x"00812d65";
		wait for Clk_period;
		Addr <=  "0101100111010";
		Trees_din <= x"ffdc2d65";
		wait for Clk_period;
		Addr <=  "0101100111011";
		Trees_din <= x"ffd82d65";
		wait for Clk_period;
		Addr <=  "0101100111100";
		Trees_din <= x"5bffb92c";
		wait for Clk_period;
		Addr <=  "0101100111101";
		Trees_din <= x"9effd820";
		wait for Clk_period;
		Addr <=  "0101100111110";
		Trees_din <= x"96ff3110";
		wait for Clk_period;
		Addr <=  "0101100111111";
		Trees_din <= x"4cfee508";
		wait for Clk_period;
		Addr <=  "0101101000000";
		Trees_din <= x"9bfef804";
		wait for Clk_period;
		Addr <=  "0101101000001";
		Trees_din <= x"00512d65";
		wait for Clk_period;
		Addr <=  "0101101000010";
		Trees_din <= x"ffa22d65";
		wait for Clk_period;
		Addr <=  "0101101000011";
		Trees_din <= x"11ffbd04";
		wait for Clk_period;
		Addr <=  "0101101000100";
		Trees_din <= x"007f2d65";
		wait for Clk_period;
		Addr <=  "0101101000101";
		Trees_din <= x"fff22d65";
		wait for Clk_period;
		Addr <=  "0101101000110";
		Trees_din <= x"5effcc08";
		wait for Clk_period;
		Addr <=  "0101101000111";
		Trees_din <= x"7efe4604";
		wait for Clk_period;
		Addr <=  "0101101001000";
		Trees_din <= x"ffc02d65";
		wait for Clk_period;
		Addr <=  "0101101001001";
		Trees_din <= x"00452d65";
		wait for Clk_period;
		Addr <=  "0101101001010";
		Trees_din <= x"d9ffe304";
		wait for Clk_period;
		Addr <=  "0101101001011";
		Trees_din <= x"000a2d65";
		wait for Clk_period;
		Addr <=  "0101101001100";
		Trees_din <= x"ff922d65";
		wait for Clk_period;
		Addr <=  "0101101001101";
		Trees_din <= x"5ffec204";
		wait for Clk_period;
		Addr <=  "0101101001110";
		Trees_din <= x"00132d65";
		wait for Clk_period;
		Addr <=  "0101101001111";
		Trees_din <= x"0700cd04";
		wait for Clk_period;
		Addr <=  "0101101010000";
		Trees_din <= x"ff7b2d65";
		wait for Clk_period;
		Addr <=  "0101101010001";
		Trees_din <= x"fff02d65";
		wait for Clk_period;
		Addr <=  "0101101010010";
		Trees_din <= x"4dfe9b08";
		wait for Clk_period;
		Addr <=  "0101101010011";
		Trees_din <= x"36ff9904";
		wait for Clk_period;
		Addr <=  "0101101010100";
		Trees_din <= x"ff6c2d65";
		wait for Clk_period;
		Addr <=  "0101101010101";
		Trees_din <= x"ffd62d65";
		wait for Clk_period;
		Addr <=  "0101101010110";
		Trees_din <= x"03ffb104";
		wait for Clk_period;
		Addr <=  "0101101010111";
		Trees_din <= x"ffd92d65";
		wait for Clk_period;
		Addr <=  "0101101011000";
		Trees_din <= x"007b2d65";
		wait for Clk_period;
		Addr <=  "0101101011001";
		Trees_din <= x"3d00295c";
		wait for Clk_period;
		Addr <=  "0101101011010";
		Trees_din <= x"97fe3a1c";
		wait for Clk_period;
		Addr <=  "0101101011011";
		Trees_din <= x"96fea908";
		wait for Clk_period;
		Addr <=  "0101101011100";
		Trees_din <= x"31ffbe04";
		wait for Clk_period;
		Addr <=  "0101101011101";
		Trees_din <= x"fff12ec1";
		wait for Clk_period;
		Addr <=  "0101101011110";
		Trees_din <= x"00692ec1";
		wait for Clk_period;
		Addr <=  "0101101011111";
		Trees_din <= x"79fe8104";
		wait for Clk_period;
		Addr <=  "0101101100000";
		Trees_din <= x"00372ec1";
		wait for Clk_period;
		Addr <=  "0101101100001";
		Trees_din <= x"8aff2d08";
		wait for Clk_period;
		Addr <=  "0101101100010";
		Trees_din <= x"b8ff1604";
		wait for Clk_period;
		Addr <=  "0101101100011";
		Trees_din <= x"005d2ec1";
		wait for Clk_period;
		Addr <=  "0101101100100";
		Trees_din <= x"ffd42ec1";
		wait for Clk_period;
		Addr <=  "0101101100101";
		Trees_din <= x"da004d04";
		wait for Clk_period;
		Addr <=  "0101101100110";
		Trees_din <= x"ff762ec1";
		wait for Clk_period;
		Addr <=  "0101101100111";
		Trees_din <= x"00142ec1";
		wait for Clk_period;
		Addr <=  "0101101101000";
		Trees_din <= x"cc004320";
		wait for Clk_period;
		Addr <=  "0101101101001";
		Trees_din <= x"61ff6710";
		wait for Clk_period;
		Addr <=  "0101101101010";
		Trees_din <= x"ddff1f08";
		wait for Clk_period;
		Addr <=  "0101101101011";
		Trees_din <= x"28ff3504";
		wait for Clk_period;
		Addr <=  "0101101101100";
		Trees_din <= x"00272ec1";
		wait for Clk_period;
		Addr <=  "0101101101101";
		Trees_din <= x"ffd12ec1";
		wait for Clk_period;
		Addr <=  "0101101101110";
		Trees_din <= x"b2ff8e04";
		wait for Clk_period;
		Addr <=  "0101101101111";
		Trees_din <= x"000c2ec1";
		wait for Clk_period;
		Addr <=  "0101101110000";
		Trees_din <= x"ffb02ec1";
		wait for Clk_period;
		Addr <=  "0101101110001";
		Trees_din <= x"7dff7508";
		wait for Clk_period;
		Addr <=  "0101101110010";
		Trees_din <= x"82001e04";
		wait for Clk_period;
		Addr <=  "0101101110011";
		Trees_din <= x"ffd42ec1";
		wait for Clk_period;
		Addr <=  "0101101110100";
		Trees_din <= x"00732ec1";
		wait for Clk_period;
		Addr <=  "0101101110101";
		Trees_din <= x"cdffe804";
		wait for Clk_period;
		Addr <=  "0101101110110";
		Trees_din <= x"002f2ec1";
		wait for Clk_period;
		Addr <=  "0101101110111";
		Trees_din <= x"fffa2ec1";
		wait for Clk_period;
		Addr <=  "0101101111000";
		Trees_din <= x"edff9910";
		wait for Clk_period;
		Addr <=  "0101101111001";
		Trees_din <= x"6bfe7308";
		wait for Clk_period;
		Addr <=  "0101101111010";
		Trees_din <= x"78ff3404";
		wait for Clk_period;
		Addr <=  "0101101111011";
		Trees_din <= x"003c2ec1";
		wait for Clk_period;
		Addr <=  "0101101111100";
		Trees_din <= x"ff9d2ec1";
		wait for Clk_period;
		Addr <=  "0101101111101";
		Trees_din <= x"aa000d04";
		wait for Clk_period;
		Addr <=  "0101101111110";
		Trees_din <= x"00772ec1";
		wait for Clk_period;
		Addr <=  "0101101111111";
		Trees_din <= x"ffbe2ec1";
		wait for Clk_period;
		Addr <=  "0101110000000";
		Trees_din <= x"02fead08";
		wait for Clk_period;
		Addr <=  "0101110000001";
		Trees_din <= x"f8001004";
		wait for Clk_period;
		Addr <=  "0101110000010";
		Trees_din <= x"005f2ec1";
		wait for Clk_period;
		Addr <=  "0101110000011";
		Trees_din <= x"ffbb2ec1";
		wait for Clk_period;
		Addr <=  "0101110000100";
		Trees_din <= x"6bfef004";
		wait for Clk_period;
		Addr <=  "0101110000101";
		Trees_din <= x"006c2ec1";
		wait for Clk_period;
		Addr <=  "0101110000110";
		Trees_din <= x"fff02ec1";
		wait for Clk_period;
		Addr <=  "0101110000111";
		Trees_din <= x"e0fe7214";
		wait for Clk_period;
		Addr <=  "0101110001000";
		Trees_din <= x"ddff6210";
		wait for Clk_period;
		Addr <=  "0101110001001";
		Trees_din <= x"a8ff0b04";
		wait for Clk_period;
		Addr <=  "0101110001010";
		Trees_din <= x"ffcd2ec1";
		wait for Clk_period;
		Addr <=  "0101110001011";
		Trees_din <= x"7cff1804";
		wait for Clk_period;
		Addr <=  "0101110001100";
		Trees_din <= x"ffff2ec1";
		wait for Clk_period;
		Addr <=  "0101110001101";
		Trees_din <= x"94ff3b04";
		wait for Clk_period;
		Addr <=  "0101110001110";
		Trees_din <= x"002c2ec1";
		wait for Clk_period;
		Addr <=  "0101110001111";
		Trees_din <= x"00a82ec1";
		wait for Clk_period;
		Addr <=  "0101110010000";
		Trees_din <= x"ffac2ec1";
		wait for Clk_period;
		Addr <=  "0101110010001";
		Trees_din <= x"7affa020";
		wait for Clk_period;
		Addr <=  "0101110010010";
		Trees_din <= x"95ff1d10";
		wait for Clk_period;
		Addr <=  "0101110010011";
		Trees_din <= x"99fede08";
		wait for Clk_period;
		Addr <=  "0101110010100";
		Trees_din <= x"cb005b04";
		wait for Clk_period;
		Addr <=  "0101110010101";
		Trees_din <= x"ff932ec1";
		wait for Clk_period;
		Addr <=  "0101110010110";
		Trees_din <= x"00662ec1";
		wait for Clk_period;
		Addr <=  "0101110010111";
		Trees_din <= x"f8006804";
		wait for Clk_period;
		Addr <=  "0101110011000";
		Trees_din <= x"00582ec1";
		wait for Clk_period;
		Addr <=  "0101110011001";
		Trees_din <= x"ffb82ec1";
		wait for Clk_period;
		Addr <=  "0101110011010";
		Trees_din <= x"6dffb008";
		wait for Clk_period;
		Addr <=  "0101110011011";
		Trees_din <= x"9effa004";
		wait for Clk_period;
		Addr <=  "0101110011100";
		Trees_din <= x"ffae2ec1";
		wait for Clk_period;
		Addr <=  "0101110011101";
		Trees_din <= x"00722ec1";
		wait for Clk_period;
		Addr <=  "0101110011110";
		Trees_din <= x"8c007c04";
		wait for Clk_period;
		Addr <=  "0101110011111";
		Trees_din <= x"ff742ec1";
		wait for Clk_period;
		Addr <=  "0101110100000";
		Trees_din <= x"001a2ec1";
		wait for Clk_period;
		Addr <=  "0101110100001";
		Trees_din <= x"56ff7d10";
		wait for Clk_period;
		Addr <=  "0101110100010";
		Trees_din <= x"94fff608";
		wait for Clk_period;
		Addr <=  "0101110100011";
		Trees_din <= x"09001b04";
		wait for Clk_period;
		Addr <=  "0101110100100";
		Trees_din <= x"ff962ec1";
		wait for Clk_period;
		Addr <=  "0101110100101";
		Trees_din <= x"00342ec1";
		wait for Clk_period;
		Addr <=  "0101110100110";
		Trees_din <= x"32fed104";
		wait for Clk_period;
		Addr <=  "0101110100111";
		Trees_din <= x"00682ec1";
		wait for Clk_period;
		Addr <=  "0101110101000";
		Trees_din <= x"ffb92ec1";
		wait for Clk_period;
		Addr <=  "0101110101001";
		Trees_din <= x"b9fed408";
		wait for Clk_period;
		Addr <=  "0101110101010";
		Trees_din <= x"5bff8204";
		wait for Clk_period;
		Addr <=  "0101110101011";
		Trees_din <= x"00192ec1";
		wait for Clk_period;
		Addr <=  "0101110101100";
		Trees_din <= x"ff822ec1";
		wait for Clk_period;
		Addr <=  "0101110101101";
		Trees_din <= x"9a006c04";
		wait for Clk_period;
		Addr <=  "0101110101110";
		Trees_din <= x"00482ec1";
		wait for Clk_period;
		Addr <=  "0101110101111";
		Trees_din <= x"ff982ec1";
		wait for Clk_period;
		Addr <=  "0101110110000";
		Trees_din <= x"6f003e74";
		wait for Clk_period;
		Addr <=  "0101110110001";
		Trees_din <= x"25007840";
		wait for Clk_period;
		Addr <=  "0101110110010";
		Trees_din <= x"9fff5920";
		wait for Clk_period;
		Addr <=  "0101110110011";
		Trees_din <= x"62ff4610";
		wait for Clk_period;
		Addr <=  "0101110110100";
		Trees_din <= x"5fffa408";
		wait for Clk_period;
		Addr <=  "0101110110101";
		Trees_din <= x"b7000b04";
		wait for Clk_period;
		Addr <=  "0101110110110";
		Trees_din <= x"00142ffd";
		wait for Clk_period;
		Addr <=  "0101110110111";
		Trees_din <= x"00502ffd";
		wait for Clk_period;
		Addr <=  "0101110111000";
		Trees_din <= x"19ff7e04";
		wait for Clk_period;
		Addr <=  "0101110111001";
		Trees_din <= x"ffa02ffd";
		wait for Clk_period;
		Addr <=  "0101110111010";
		Trees_din <= x"00352ffd";
		wait for Clk_period;
		Addr <=  "0101110111011";
		Trees_din <= x"f9ff2f08";
		wait for Clk_period;
		Addr <=  "0101110111100";
		Trees_din <= x"9bffa304";
		wait for Clk_period;
		Addr <=  "0101110111101";
		Trees_din <= x"fff92ffd";
		wait for Clk_period;
		Addr <=  "0101110111110";
		Trees_din <= x"005a2ffd";
		wait for Clk_period;
		Addr <=  "0101110111111";
		Trees_din <= x"2a015804";
		wait for Clk_period;
		Addr <=  "0101111000000";
		Trees_din <= x"ffb82ffd";
		wait for Clk_period;
		Addr <=  "0101111000001";
		Trees_din <= x"00402ffd";
		wait for Clk_period;
		Addr <=  "0101111000010";
		Trees_din <= x"55ffd310";
		wait for Clk_period;
		Addr <=  "0101111000011";
		Trees_din <= x"9bff9108";
		wait for Clk_period;
		Addr <=  "0101111000100";
		Trees_din <= x"8eff8e04";
		wait for Clk_period;
		Addr <=  "0101111000101";
		Trees_din <= x"ffaf2ffd";
		wait for Clk_period;
		Addr <=  "0101111000110";
		Trees_din <= x"00312ffd";
		wait for Clk_period;
		Addr <=  "0101111000111";
		Trees_din <= x"83fea504";
		wait for Clk_period;
		Addr <=  "0101111001000";
		Trees_din <= x"003c2ffd";
		wait for Clk_period;
		Addr <=  "0101111001001";
		Trees_din <= x"ff892ffd";
		wait for Clk_period;
		Addr <=  "0101111001010";
		Trees_din <= x"5fff2308";
		wait for Clk_period;
		Addr <=  "0101111001011";
		Trees_din <= x"d6006204";
		wait for Clk_period;
		Addr <=  "0101111001100";
		Trees_din <= x"ff932ffd";
		wait for Clk_period;
		Addr <=  "0101111001101";
		Trees_din <= x"ffe02ffd";
		wait for Clk_period;
		Addr <=  "0101111001110";
		Trees_din <= x"c7ff8a04";
		wait for Clk_period;
		Addr <=  "0101111001111";
		Trees_din <= x"fff72ffd";
		wait for Clk_period;
		Addr <=  "0101111010000";
		Trees_din <= x"ff772ffd";
		wait for Clk_period;
		Addr <=  "0101111010001";
		Trees_din <= x"fdff9b20";
		wait for Clk_period;
		Addr <=  "0101111010010";
		Trees_din <= x"34ffe410";
		wait for Clk_period;
		Addr <=  "0101111010011";
		Trees_din <= x"77ff3d08";
		wait for Clk_period;
		Addr <=  "0101111010100";
		Trees_din <= x"7efece04";
		wait for Clk_period;
		Addr <=  "0101111010101";
		Trees_din <= x"fff92ffd";
		wait for Clk_period;
		Addr <=  "0101111010110";
		Trees_din <= x"ff702ffd";
		wait for Clk_period;
		Addr <=  "0101111010111";
		Trees_din <= x"f3fe8904";
		wait for Clk_period;
		Addr <=  "0101111011000";
		Trees_din <= x"ffbc2ffd";
		wait for Clk_period;
		Addr <=  "0101111011001";
		Trees_din <= x"006b2ffd";
		wait for Clk_period;
		Addr <=  "0101111011010";
		Trees_din <= x"89fffd08";
		wait for Clk_period;
		Addr <=  "0101111011011";
		Trees_din <= x"bcfefb04";
		wait for Clk_period;
		Addr <=  "0101111011100";
		Trees_din <= x"00832ffd";
		wait for Clk_period;
		Addr <=  "0101111011101";
		Trees_din <= x"002b2ffd";
		wait for Clk_period;
		Addr <=  "0101111011110";
		Trees_din <= x"72001604";
		wait for Clk_period;
		Addr <=  "0101111011111";
		Trees_din <= x"004c2ffd";
		wait for Clk_period;
		Addr <=  "0101111100000";
		Trees_din <= x"ffe62ffd";
		wait for Clk_period;
		Addr <=  "0101111100001";
		Trees_din <= x"a2002e10";
		wait for Clk_period;
		Addr <=  "0101111100010";
		Trees_din <= x"eaff4708";
		wait for Clk_period;
		Addr <=  "0101111100011";
		Trees_din <= x"21ff9904";
		wait for Clk_period;
		Addr <=  "0101111100100";
		Trees_din <= x"00522ffd";
		wait for Clk_period;
		Addr <=  "0101111100101";
		Trees_din <= x"ffd62ffd";
		wait for Clk_period;
		Addr <=  "0101111100110";
		Trees_din <= x"48ff9504";
		wait for Clk_period;
		Addr <=  "0101111100111";
		Trees_din <= x"fffe2ffd";
		wait for Clk_period;
		Addr <=  "0101111101000";
		Trees_din <= x"ff8f2ffd";
		wait for Clk_period;
		Addr <=  "0101111101001";
		Trees_din <= x"009a2ffd";
		wait for Clk_period;
		Addr <=  "0101111101010";
		Trees_din <= x"f6fec10c";
		wait for Clk_period;
		Addr <=  "0101111101011";
		Trees_din <= x"37ffe208";
		wait for Clk_period;
		Addr <=  "0101111101100";
		Trees_din <= x"6f005e04";
		wait for Clk_period;
		Addr <=  "0101111101101";
		Trees_din <= x"ffcc2ffd";
		wait for Clk_period;
		Addr <=  "0101111101110";
		Trees_din <= x"00522ffd";
		wait for Clk_period;
		Addr <=  "0101111101111";
		Trees_din <= x"ff902ffd";
		wait for Clk_period;
		Addr <=  "0101111110000";
		Trees_din <= x"7aff5c0c";
		wait for Clk_period;
		Addr <=  "0101111110001";
		Trees_din <= x"90ff5808";
		wait for Clk_period;
		Addr <=  "0101111110010";
		Trees_din <= x"f202e204";
		wait for Clk_period;
		Addr <=  "0101111110011";
		Trees_din <= x"fff62ffd";
		wait for Clk_period;
		Addr <=  "0101111110100";
		Trees_din <= x"00742ffd";
		wait for Clk_period;
		Addr <=  "0101111110101";
		Trees_din <= x"ffa12ffd";
		wait for Clk_period;
		Addr <=  "0101111110110";
		Trees_din <= x"bfff6108";
		wait for Clk_period;
		Addr <=  "0101111110111";
		Trees_din <= x"53ff8704";
		wait for Clk_period;
		Addr <=  "0101111111000";
		Trees_din <= x"ff9f2ffd";
		wait for Clk_period;
		Addr <=  "0101111111001";
		Trees_din <= x"00542ffd";
		wait for Clk_period;
		Addr <=  "0101111111010";
		Trees_din <= x"aafee904";
		wait for Clk_period;
		Addr <=  "0101111111011";
		Trees_din <= x"ffe52ffd";
		wait for Clk_period;
		Addr <=  "0101111111100";
		Trees_din <= x"9eff6f04";
		wait for Clk_period;
		Addr <=  "0101111111101";
		Trees_din <= x"00402ffd";
		wait for Clk_period;
		Addr <=  "0101111111110";
		Trees_din <= x"00b12ffd";
		wait for Clk_period;
		Addr <=  "0101111111111";
		Trees_din <= x"3cff7e58";
		wait for Clk_period;
		Addr <=  "0110000000000";
		Trees_din <= x"8ffe011c";
		wait for Clk_period;
		Addr <=  "0110000000001";
		Trees_din <= x"b0ff150c";
		wait for Clk_period;
		Addr <=  "0110000000010";
		Trees_din <= x"91ff5608";
		wait for Clk_period;
		Addr <=  "0110000000011";
		Trees_din <= x"34001304";
		wait for Clk_period;
		Addr <=  "0110000000100";
		Trees_din <= x"008430f1";
		wait for Clk_period;
		Addr <=  "0110000000101";
		Trees_din <= x"ffe130f1";
		wait for Clk_period;
		Addr <=  "0110000000110";
		Trees_din <= x"ffad30f1";
		wait for Clk_period;
		Addr <=  "0110000000111";
		Trees_din <= x"09fec804";
		wait for Clk_period;
		Addr <=  "0110000001000";
		Trees_din <= x"005830f1";
		wait for Clk_period;
		Addr <=  "0110000001001";
		Trees_din <= x"cd007208";
		wait for Clk_period;
		Addr <=  "0110000001010";
		Trees_din <= x"2aff1a04";
		wait for Clk_period;
		Addr <=  "0110000001011";
		Trees_din <= x"fffe30f1";
		wait for Clk_period;
		Addr <=  "0110000001100";
		Trees_din <= x"ff7030f1";
		wait for Clk_period;
		Addr <=  "0110000001101";
		Trees_din <= x"003930f1";
		wait for Clk_period;
		Addr <=  "0110000001110";
		Trees_din <= x"33fec21c";
		wait for Clk_period;
		Addr <=  "0110000001111";
		Trees_din <= x"24ffc910";
		wait for Clk_period;
		Addr <=  "0110000010000";
		Trees_din <= x"11ffb708";
		wait for Clk_period;
		Addr <=  "0110000010001";
		Trees_din <= x"cf005404";
		wait for Clk_period;
		Addr <=  "0110000010010";
		Trees_din <= x"002b30f1";
		wait for Clk_period;
		Addr <=  "0110000010011";
		Trees_din <= x"008030f1";
		wait for Clk_period;
		Addr <=  "0110000010100";
		Trees_din <= x"cafea804";
		wait for Clk_period;
		Addr <=  "0110000010101";
		Trees_din <= x"ffa230f1";
		wait for Clk_period;
		Addr <=  "0110000010110";
		Trees_din <= x"006230f1";
		wait for Clk_period;
		Addr <=  "0110000010111";
		Trees_din <= x"4fff1404";
		wait for Clk_period;
		Addr <=  "0110000011000";
		Trees_din <= x"ff9330f1";
		wait for Clk_period;
		Addr <=  "0110000011001";
		Trees_din <= x"7cffc504";
		wait for Clk_period;
		Addr <=  "0110000011010";
		Trees_din <= x"003230f1";
		wait for Clk_period;
		Addr <=  "0110000011011";
		Trees_din <= x"ffcf30f1";
		wait for Clk_period;
		Addr <=  "0110000011100";
		Trees_din <= x"5d001110";
		wait for Clk_period;
		Addr <=  "0110000011101";
		Trees_din <= x"3cff5f08";
		wait for Clk_period;
		Addr <=  "0110000011110";
		Trees_din <= x"a1ffab04";
		wait for Clk_period;
		Addr <=  "0110000011111";
		Trees_din <= x"000830f1";
		wait for Clk_period;
		Addr <=  "0110000100000";
		Trees_din <= x"ffd530f1";
		wait for Clk_period;
		Addr <=  "0110000100001";
		Trees_din <= x"e1ffd404";
		wait for Clk_period;
		Addr <=  "0110000100010";
		Trees_din <= x"006130f1";
		wait for Clk_period;
		Addr <=  "0110000100011";
		Trees_din <= x"fff130f1";
		wait for Clk_period;
		Addr <=  "0110000100100";
		Trees_din <= x"f8fffe08";
		wait for Clk_period;
		Addr <=  "0110000100101";
		Trees_din <= x"bcfedc04";
		wait for Clk_period;
		Addr <=  "0110000100110";
		Trees_din <= x"008730f1";
		wait for Clk_period;
		Addr <=  "0110000100111";
		Trees_din <= x"ffdd30f1";
		wait for Clk_period;
		Addr <=  "0110000101000";
		Trees_din <= x"2bff7e04";
		wait for Clk_period;
		Addr <=  "0110000101001";
		Trees_din <= x"001230f1";
		wait for Clk_period;
		Addr <=  "0110000101010";
		Trees_din <= x"ffa930f1";
		wait for Clk_period;
		Addr <=  "0110000101011";
		Trees_din <= x"47001c0c";
		wait for Clk_period;
		Addr <=  "0110000101100";
		Trees_din <= x"f7fef904";
		wait for Clk_period;
		Addr <=  "0110000101101";
		Trees_din <= x"001730f1";
		wait for Clk_period;
		Addr <=  "0110000101110";
		Trees_din <= x"41fe9604";
		wait for Clk_period;
		Addr <=  "0110000101111";
		Trees_din <= x"ffea30f1";
		wait for Clk_period;
		Addr <=  "0110000110000";
		Trees_din <= x"ff6d30f1";
		wait for Clk_period;
		Addr <=  "0110000110001";
		Trees_din <= x"8fff210c";
		wait for Clk_period;
		Addr <=  "0110000110010";
		Trees_din <= x"c0ff5404";
		wait for Clk_period;
		Addr <=  "0110000110011";
		Trees_din <= x"ffbe30f1";
		wait for Clk_period;
		Addr <=  "0110000110100";
		Trees_din <= x"35ff0e04";
		wait for Clk_period;
		Addr <=  "0110000110101";
		Trees_din <= x"008c30f1";
		wait for Clk_period;
		Addr <=  "0110000110110";
		Trees_din <= x"ffff30f1";
		wait for Clk_period;
		Addr <=  "0110000110111";
		Trees_din <= x"63ff4e04";
		wait for Clk_period;
		Addr <=  "0110000111000";
		Trees_din <= x"003630f1";
		wait for Clk_period;
		Addr <=  "0110000111001";
		Trees_din <= x"50ff4904";
		wait for Clk_period;
		Addr <=  "0110000111010";
		Trees_din <= x"ffdf30f1";
		wait for Clk_period;
		Addr <=  "0110000111011";
		Trees_din <= x"ff8530f1";
		wait for Clk_period;
		Addr <=  "0110000111100";
		Trees_din <= x"44005368";
		wait for Clk_period;
		Addr <=  "0110000111101";
		Trees_din <= x"60ffcd40";
		wait for Clk_period;
		Addr <=  "0110000111110";
		Trees_din <= x"2dff1320";
		wait for Clk_period;
		Addr <=  "0110000111111";
		Trees_din <= x"71fff110";
		wait for Clk_period;
		Addr <=  "0110001000000";
		Trees_din <= x"9cfeec08";
		wait for Clk_period;
		Addr <=  "0110001000001";
		Trees_din <= x"3aff9104";
		wait for Clk_period;
		Addr <=  "0110001000010";
		Trees_din <= x"004a321d";
		wait for Clk_period;
		Addr <=  "0110001000011";
		Trees_din <= x"ffe4321d";
		wait for Clk_period;
		Addr <=  "0110001000100";
		Trees_din <= x"55ff9304";
		wait for Clk_period;
		Addr <=  "0110001000101";
		Trees_din <= x"0023321d";
		wait for Clk_period;
		Addr <=  "0110001000110";
		Trees_din <= x"ffd4321d";
		wait for Clk_period;
		Addr <=  "0110001000111";
		Trees_din <= x"c3002608";
		wait for Clk_period;
		Addr <=  "0110001001000";
		Trees_din <= x"47003a04";
		wait for Clk_period;
		Addr <=  "0110001001001";
		Trees_din <= x"ffac321d";
		wait for Clk_period;
		Addr <=  "0110001001010";
		Trees_din <= x"0033321d";
		wait for Clk_period;
		Addr <=  "0110001001011";
		Trees_din <= x"d5ffae04";
		wait for Clk_period;
		Addr <=  "0110001001100";
		Trees_din <= x"0002321d";
		wait for Clk_period;
		Addr <=  "0110001001101";
		Trees_din <= x"0085321d";
		wait for Clk_period;
		Addr <=  "0110001001110";
		Trees_din <= x"cbffed10";
		wait for Clk_period;
		Addr <=  "0110001001111";
		Trees_din <= x"01ff4308";
		wait for Clk_period;
		Addr <=  "0110001010000";
		Trees_din <= x"c6ffad04";
		wait for Clk_period;
		Addr <=  "0110001010001";
		Trees_din <= x"0032321d";
		wait for Clk_period;
		Addr <=  "0110001010010";
		Trees_din <= x"ffdd321d";
		wait for Clk_period;
		Addr <=  "0110001010011";
		Trees_din <= x"59ff3f04";
		wait for Clk_period;
		Addr <=  "0110001010100";
		Trees_din <= x"0028321d";
		wait for Clk_period;
		Addr <=  "0110001010101";
		Trees_din <= x"ff99321d";
		wait for Clk_period;
		Addr <=  "0110001010110";
		Trees_din <= x"cdffd008";
		wait for Clk_period;
		Addr <=  "0110001010111";
		Trees_din <= x"6bfef304";
		wait for Clk_period;
		Addr <=  "0110001011000";
		Trees_din <= x"002e321d";
		wait for Clk_period;
		Addr <=  "0110001011001";
		Trees_din <= x"ff9f321d";
		wait for Clk_period;
		Addr <=  "0110001011010";
		Trees_din <= x"8bff8f04";
		wait for Clk_period;
		Addr <=  "0110001011011";
		Trees_din <= x"0040321d";
		wait for Clk_period;
		Addr <=  "0110001011100";
		Trees_din <= x"ff91321d";
		wait for Clk_period;
		Addr <=  "0110001011101";
		Trees_din <= x"0d001f14";
		wait for Clk_period;
		Addr <=  "0110001011110";
		Trees_din <= x"95fff210";
		wait for Clk_period;
		Addr <=  "0110001011111";
		Trees_din <= x"56ff7d08";
		wait for Clk_period;
		Addr <=  "0110001100000";
		Trees_din <= x"3bff7c04";
		wait for Clk_period;
		Addr <=  "0110001100001";
		Trees_din <= x"ffee321d";
		wait for Clk_period;
		Addr <=  "0110001100010";
		Trees_din <= x"0044321d";
		wait for Clk_period;
		Addr <=  "0110001100011";
		Trees_din <= x"8ffe5204";
		wait for Clk_period;
		Addr <=  "0110001100100";
		Trees_din <= x"ffb2321d";
		wait for Clk_period;
		Addr <=  "0110001100101";
		Trees_din <= x"0056321d";
		wait for Clk_period;
		Addr <=  "0110001100110";
		Trees_din <= x"ff8a321d";
		wait for Clk_period;
		Addr <=  "0110001100111";
		Trees_din <= x"be00340c";
		wait for Clk_period;
		Addr <=  "0110001101000";
		Trees_din <= x"a5ff5f08";
		wait for Clk_period;
		Addr <=  "0110001101001";
		Trees_din <= x"95feb404";
		wait for Clk_period;
		Addr <=  "0110001101010";
		Trees_din <= x"ffdb321d";
		wait for Clk_period;
		Addr <=  "0110001101011";
		Trees_din <= x"ff77321d";
		wait for Clk_period;
		Addr <=  "0110001101100";
		Trees_din <= x"001c321d";
		wait for Clk_period;
		Addr <=  "0110001101101";
		Trees_din <= x"27ffa604";
		wait for Clk_period;
		Addr <=  "0110001101110";
		Trees_din <= x"006e321d";
		wait for Clk_period;
		Addr <=  "0110001101111";
		Trees_din <= x"ffc3321d";
		wait for Clk_period;
		Addr <=  "0110001110000";
		Trees_din <= x"eaffe924";
		wait for Clk_period;
		Addr <=  "0110001110001";
		Trees_din <= x"30007120";
		wait for Clk_period;
		Addr <=  "0110001110010";
		Trees_din <= x"96ff2a10";
		wait for Clk_period;
		Addr <=  "0110001110011";
		Trees_din <= x"4cfee508";
		wait for Clk_period;
		Addr <=  "0110001110100";
		Trees_din <= x"44008c04";
		wait for Clk_period;
		Addr <=  "0110001110101";
		Trees_din <= x"ff9e321d";
		wait for Clk_period;
		Addr <=  "0110001110110";
		Trees_din <= x"0043321d";
		wait for Clk_period;
		Addr <=  "0110001110111";
		Trees_din <= x"e7fee404";
		wait for Clk_period;
		Addr <=  "0110001111000";
		Trees_din <= x"ffc7321d";
		wait for Clk_period;
		Addr <=  "0110001111001";
		Trees_din <= x"0071321d";
		wait for Clk_period;
		Addr <=  "0110001111010";
		Trees_din <= x"5effcc08";
		wait for Clk_period;
		Addr <=  "0110001111011";
		Trees_din <= x"faff7004";
		wait for Clk_period;
		Addr <=  "0110001111100";
		Trees_din <= x"0003321d";
		wait for Clk_period;
		Addr <=  "0110001111101";
		Trees_din <= x"0064321d";
		wait for Clk_period;
		Addr <=  "0110001111110";
		Trees_din <= x"b3fee704";
		wait for Clk_period;
		Addr <=  "0110001111111";
		Trees_din <= x"0042321d";
		wait for Clk_period;
		Addr <=  "0110010000000";
		Trees_din <= x"ffc7321d";
		wait for Clk_period;
		Addr <=  "0110010000001";
		Trees_din <= x"ff8f321d";
		wait for Clk_period;
		Addr <=  "0110010000010";
		Trees_din <= x"ba000108";
		wait for Clk_period;
		Addr <=  "0110010000011";
		Trees_din <= x"1eff3404";
		wait for Clk_period;
		Addr <=  "0110010000100";
		Trees_din <= x"ffe4321d";
		wait for Clk_period;
		Addr <=  "0110010000101";
		Trees_din <= x"ff82321d";
		wait for Clk_period;
		Addr <=  "0110010000110";
		Trees_din <= x"0021321d";
		wait for Clk_period;
		Addr <=  "0110010000111";
		Trees_din <= x"f3fee544";
		wait for Clk_period;
		Addr <=  "0110010001000";
		Trees_din <= x"a1fff83c";
		wait for Clk_period;
		Addr <=  "0110010001001";
		Trees_din <= x"e3ff1820";
		wait for Clk_period;
		Addr <=  "0110010001010";
		Trees_din <= x"45ff4710";
		wait for Clk_period;
		Addr <=  "0110010001011";
		Trees_din <= x"8800ec08";
		wait for Clk_period;
		Addr <=  "0110010001100";
		Trees_din <= x"c1fe7204";
		wait for Clk_period;
		Addr <=  "0110010001101";
		Trees_din <= x"fff53349";
		wait for Clk_period;
		Addr <=  "0110010001110";
		Trees_din <= x"00283349";
		wait for Clk_period;
		Addr <=  "0110010001111";
		Trees_din <= x"93ffe104";
		wait for Clk_period;
		Addr <=  "0110010010000";
		Trees_din <= x"ff883349";
		wait for Clk_period;
		Addr <=  "0110010010001";
		Trees_din <= x"00143349";
		wait for Clk_period;
		Addr <=  "0110010010010";
		Trees_din <= x"dbffc808";
		wait for Clk_period;
		Addr <=  "0110010010011";
		Trees_din <= x"66001e04";
		wait for Clk_period;
		Addr <=  "0110010010100";
		Trees_din <= x"ff783349";
		wait for Clk_period;
		Addr <=  "0110010010101";
		Trees_din <= x"00403349";
		wait for Clk_period;
		Addr <=  "0110010010110";
		Trees_din <= x"02ff0c04";
		wait for Clk_period;
		Addr <=  "0110010010111";
		Trees_din <= x"00213349";
		wait for Clk_period;
		Addr <=  "0110010011000";
		Trees_din <= x"ffaf3349";
		wait for Clk_period;
		Addr <=  "0110010011001";
		Trees_din <= x"c5ff5d10";
		wait for Clk_period;
		Addr <=  "0110010011010";
		Trees_din <= x"60fff108";
		wait for Clk_period;
		Addr <=  "0110010011011";
		Trees_din <= x"0bff2804";
		wait for Clk_period;
		Addr <=  "0110010011100";
		Trees_din <= x"00343349";
		wait for Clk_period;
		Addr <=  "0110010011101";
		Trees_din <= x"ff813349";
		wait for Clk_period;
		Addr <=  "0110010011110";
		Trees_din <= x"3eff7804";
		wait for Clk_period;
		Addr <=  "0110010011111";
		Trees_din <= x"ffe63349";
		wait for Clk_period;
		Addr <=  "0110010100000";
		Trees_din <= x"00763349";
		wait for Clk_period;
		Addr <=  "0110010100001";
		Trees_din <= x"5dfff408";
		wait for Clk_period;
		Addr <=  "0110010100010";
		Trees_din <= x"d3fef504";
		wait for Clk_period;
		Addr <=  "0110010100011";
		Trees_din <= x"fff93349";
		wait for Clk_period;
		Addr <=  "0110010100100";
		Trees_din <= x"00933349";
		wait for Clk_period;
		Addr <=  "0110010100101";
		Trees_din <= x"ffad3349";
		wait for Clk_period;
		Addr <=  "0110010100110";
		Trees_din <= x"52ff0504";
		wait for Clk_period;
		Addr <=  "0110010100111";
		Trees_din <= x"001f3349";
		wait for Clk_period;
		Addr <=  "0110010101000";
		Trees_din <= x"ff7f3349";
		wait for Clk_period;
		Addr <=  "0110010101001";
		Trees_din <= x"00ffdc40";
		wait for Clk_period;
		Addr <=  "0110010101010";
		Trees_din <= x"05005f20";
		wait for Clk_period;
		Addr <=  "0110010101011";
		Trees_din <= x"faffc510";
		wait for Clk_period;
		Addr <=  "0110010101100";
		Trees_din <= x"0affc408";
		wait for Clk_period;
		Addr <=  "0110010101101";
		Trees_din <= x"bdff9c04";
		wait for Clk_period;
		Addr <=  "0110010101110";
		Trees_din <= x"00483349";
		wait for Clk_period;
		Addr <=  "0110010101111";
		Trees_din <= x"ffd63349";
		wait for Clk_period;
		Addr <=  "0110010110000";
		Trees_din <= x"97ff6e04";
		wait for Clk_period;
		Addr <=  "0110010110001";
		Trees_din <= x"ffb43349";
		wait for Clk_period;
		Addr <=  "0110010110010";
		Trees_din <= x"00053349";
		wait for Clk_period;
		Addr <=  "0110010110011";
		Trees_din <= x"5dffb008";
		wait for Clk_period;
		Addr <=  "0110010110100";
		Trees_din <= x"27ff8004";
		wait for Clk_period;
		Addr <=  "0110010110101";
		Trees_din <= x"ffc83349";
		wait for Clk_period;
		Addr <=  "0110010110110";
		Trees_din <= x"007e3349";
		wait for Clk_period;
		Addr <=  "0110010110111";
		Trees_din <= x"a0ff4404";
		wait for Clk_period;
		Addr <=  "0110010111000";
		Trees_din <= x"ffa23349";
		wait for Clk_period;
		Addr <=  "0110010111001";
		Trees_din <= x"00373349";
		wait for Clk_period;
		Addr <=  "0110010111010";
		Trees_din <= x"52ff8010";
		wait for Clk_period;
		Addr <=  "0110010111011";
		Trees_din <= x"0bff7408";
		wait for Clk_period;
		Addr <=  "0110010111100";
		Trees_din <= x"29ff9404";
		wait for Clk_period;
		Addr <=  "0110010111101";
		Trees_din <= x"ff993349";
		wait for Clk_period;
		Addr <=  "0110010111110";
		Trees_din <= x"00203349";
		wait for Clk_period;
		Addr <=  "0110010111111";
		Trees_din <= x"58feea04";
		wait for Clk_period;
		Addr <=  "0110011000000";
		Trees_din <= x"00433349";
		wait for Clk_period;
		Addr <=  "0110011000001";
		Trees_din <= x"00073349";
		wait for Clk_period;
		Addr <=  "0110011000010";
		Trees_din <= x"d7008b08";
		wait for Clk_period;
		Addr <=  "0110011000011";
		Trees_din <= x"f3ffce04";
		wait for Clk_period;
		Addr <=  "0110011000100";
		Trees_din <= x"ff883349";
		wait for Clk_period;
		Addr <=  "0110011000101";
		Trees_din <= x"001c3349";
		wait for Clk_period;
		Addr <=  "0110011000110";
		Trees_din <= x"35fed604";
		wait for Clk_period;
		Addr <=  "0110011000111";
		Trees_din <= x"004a3349";
		wait for Clk_period;
		Addr <=  "0110011001000";
		Trees_din <= x"ffc63349";
		wait for Clk_period;
		Addr <=  "0110011001001";
		Trees_din <= x"effeef08";
		wait for Clk_period;
		Addr <=  "0110011001010";
		Trees_din <= x"92ff2704";
		wait for Clk_period;
		Addr <=  "0110011001011";
		Trees_din <= x"ffc13349";
		wait for Clk_period;
		Addr <=  "0110011001100";
		Trees_din <= x"00543349";
		wait for Clk_period;
		Addr <=  "0110011001101";
		Trees_din <= x"b7000f08";
		wait for Clk_period;
		Addr <=  "0110011001110";
		Trees_din <= x"64ff9804";
		wait for Clk_period;
		Addr <=  "0110011001111";
		Trees_din <= x"ff6e3349";
		wait for Clk_period;
		Addr <=  "0110011010000";
		Trees_din <= x"ffde3349";
		wait for Clk_period;
		Addr <=  "0110011010001";
		Trees_din <= x"00183349";
		wait for Clk_period;
		Addr <=  "0110011010010";
		Trees_din <= x"2eff354c";
		wait for Clk_period;
		Addr <=  "0110011010011";
		Trees_din <= x"e6ffc12c";
		wait for Clk_period;
		Addr <=  "0110011010100";
		Trees_din <= x"8aff8414";
		wait for Clk_period;
		Addr <=  "0110011010101";
		Trees_din <= x"31ff8108";
		wait for Clk_period;
		Addr <=  "0110011010110";
		Trees_din <= x"7efe6f04";
		wait for Clk_period;
		Addr <=  "0110011010111";
		Trees_din <= x"002c34b5";
		wait for Clk_period;
		Addr <=  "0110011011000";
		Trees_din <= x"ff9534b5";
		wait for Clk_period;
		Addr <=  "0110011011001";
		Trees_din <= x"50ff4604";
		wait for Clk_period;
		Addr <=  "0110011011010";
		Trees_din <= x"ffe234b5";
		wait for Clk_period;
		Addr <=  "0110011011011";
		Trees_din <= x"2cffd104";
		wait for Clk_period;
		Addr <=  "0110011011100";
		Trees_din <= x"009734b5";
		wait for Clk_period;
		Addr <=  "0110011011101";
		Trees_din <= x"002c34b5";
		wait for Clk_period;
		Addr <=  "0110011011110";
		Trees_din <= x"6bfee510";
		wait for Clk_period;
		Addr <=  "0110011011111";
		Trees_din <= x"08008908";
		wait for Clk_period;
		Addr <=  "0110011100000";
		Trees_din <= x"bfff6704";
		wait for Clk_period;
		Addr <=  "0110011100001";
		Trees_din <= x"001934b5";
		wait for Clk_period;
		Addr <=  "0110011100010";
		Trees_din <= x"ff9c34b5";
		wait for Clk_period;
		Addr <=  "0110011100011";
		Trees_din <= x"f4fef504";
		wait for Clk_period;
		Addr <=  "0110011100100";
		Trees_din <= x"006234b5";
		wait for Clk_period;
		Addr <=  "0110011100101";
		Trees_din <= x"ffce34b5";
		wait for Clk_period;
		Addr <=  "0110011100110";
		Trees_din <= x"dbff9604";
		wait for Clk_period;
		Addr <=  "0110011100111";
		Trees_din <= x"fff534b5";
		wait for Clk_period;
		Addr <=  "0110011101000";
		Trees_din <= x"ff7734b5";
		wait for Clk_period;
		Addr <=  "0110011101001";
		Trees_din <= x"05000208";
		wait for Clk_period;
		Addr <=  "0110011101010";
		Trees_din <= x"adffdb04";
		wait for Clk_period;
		Addr <=  "0110011101011";
		Trees_din <= x"ff9f34b5";
		wait for Clk_period;
		Addr <=  "0110011101100";
		Trees_din <= x"003c34b5";
		wait for Clk_period;
		Addr <=  "0110011101101";
		Trees_din <= x"ec001d0c";
		wait for Clk_period;
		Addr <=  "0110011101110";
		Trees_din <= x"65000c08";
		wait for Clk_period;
		Addr <=  "0110011101111";
		Trees_din <= x"3cff8404";
		wait for Clk_period;
		Addr <=  "0110011110000";
		Trees_din <= x"007834b5";
		wait for Clk_period;
		Addr <=  "0110011110001";
		Trees_din <= x"ffd734b5";
		wait for Clk_period;
		Addr <=  "0110011110010";
		Trees_din <= x"ffc434b5";
		wait for Clk_period;
		Addr <=  "0110011110011";
		Trees_din <= x"03ffd604";
		wait for Clk_period;
		Addr <=  "0110011110100";
		Trees_din <= x"ff9934b5";
		wait for Clk_period;
		Addr <=  "0110011110101";
		Trees_din <= x"81ffbc04";
		wait for Clk_period;
		Addr <=  "0110011110110";
		Trees_din <= x"007234b5";
		wait for Clk_period;
		Addr <=  "0110011110111";
		Trees_din <= x"ffe334b5";
		wait for Clk_period;
		Addr <=  "0110011111000";
		Trees_din <= x"cffffc34";
		wait for Clk_period;
		Addr <=  "0110011111001";
		Trees_din <= x"40fffe14";
		wait for Clk_period;
		Addr <=  "0110011111010";
		Trees_din <= x"89fee304";
		wait for Clk_period;
		Addr <=  "0110011111011";
		Trees_din <= x"005a34b5";
		wait for Clk_period;
		Addr <=  "0110011111100";
		Trees_din <= x"6effe008";
		wait for Clk_period;
		Addr <=  "0110011111101";
		Trees_din <= x"15ff6504";
		wait for Clk_period;
		Addr <=  "0110011111110";
		Trees_din <= x"ffa434b5";
		wait for Clk_period;
		Addr <=  "0110011111111";
		Trees_din <= x"003734b5";
		wait for Clk_period;
		Addr <=  "0110100000000";
		Trees_din <= x"8c008404";
		wait for Clk_period;
		Addr <=  "0110100000001";
		Trees_din <= x"ff7c34b5";
		wait for Clk_period;
		Addr <=  "0110100000010";
		Trees_din <= x"000434b5";
		wait for Clk_period;
		Addr <=  "0110100000011";
		Trees_din <= x"5bff8e10";
		wait for Clk_period;
		Addr <=  "0110100000100";
		Trees_din <= x"9bfef008";
		wait for Clk_period;
		Addr <=  "0110100000101";
		Trees_din <= x"fcff3f04";
		wait for Clk_period;
		Addr <=  "0110100000110";
		Trees_din <= x"006034b5";
		wait for Clk_period;
		Addr <=  "0110100000111";
		Trees_din <= x"ffe034b5";
		wait for Clk_period;
		Addr <=  "0110100001000";
		Trees_din <= x"9dfffc04";
		wait for Clk_period;
		Addr <=  "0110100001001";
		Trees_din <= x"ffdc34b5";
		wait for Clk_period;
		Addr <=  "0110100001010";
		Trees_din <= x"004134b5";
		wait for Clk_period;
		Addr <=  "0110100001011";
		Trees_din <= x"b5fe7308";
		wait for Clk_period;
		Addr <=  "0110100001100";
		Trees_din <= x"23ff5804";
		wait for Clk_period;
		Addr <=  "0110100001101";
		Trees_din <= x"ffa734b5";
		wait for Clk_period;
		Addr <=  "0110100001110";
		Trees_din <= x"004134b5";
		wait for Clk_period;
		Addr <=  "0110100001111";
		Trees_din <= x"2ffef004";
		wait for Clk_period;
		Addr <=  "0110100010000";
		Trees_din <= x"002b34b5";
		wait for Clk_period;
		Addr <=  "0110100010001";
		Trees_din <= x"ff9834b5";
		wait for Clk_period;
		Addr <=  "0110100010010";
		Trees_din <= x"7cff8420";
		wait for Clk_period;
		Addr <=  "0110100010011";
		Trees_din <= x"d6007c10";
		wait for Clk_period;
		Addr <=  "0110100010100";
		Trees_din <= x"1afe7f08";
		wait for Clk_period;
		Addr <=  "0110100010101";
		Trees_din <= x"98fe6604";
		wait for Clk_period;
		Addr <=  "0110100010110";
		Trees_din <= x"005334b5";
		wait for Clk_period;
		Addr <=  "0110100010111";
		Trees_din <= x"ffab34b5";
		wait for Clk_period;
		Addr <=  "0110100011000";
		Trees_din <= x"9affb104";
		wait for Clk_period;
		Addr <=  "0110100011001";
		Trees_din <= x"004234b5";
		wait for Clk_period;
		Addr <=  "0110100011010";
		Trees_din <= x"ffff34b5";
		wait for Clk_period;
		Addr <=  "0110100011011";
		Trees_din <= x"30fff908";
		wait for Clk_period;
		Addr <=  "0110100011100";
		Trees_din <= x"8ffe3d04";
		wait for Clk_period;
		Addr <=  "0110100011101";
		Trees_din <= x"ffc334b5";
		wait for Clk_period;
		Addr <=  "0110100011110";
		Trees_din <= x"006034b5";
		wait for Clk_period;
		Addr <=  "0110100011111";
		Trees_din <= x"73ffe704";
		wait for Clk_period;
		Addr <=  "0110100100000";
		Trees_din <= x"ffb034b5";
		wait for Clk_period;
		Addr <=  "0110100100001";
		Trees_din <= x"003b34b5";
		wait for Clk_period;
		Addr <=  "0110100100010";
		Trees_din <= x"3b003510";
		wait for Clk_period;
		Addr <=  "0110100100011";
		Trees_din <= x"75ff8e08";
		wait for Clk_period;
		Addr <=  "0110100100100";
		Trees_din <= x"40006904";
		wait for Clk_period;
		Addr <=  "0110100100101";
		Trees_din <= x"ffa034b5";
		wait for Clk_period;
		Addr <=  "0110100100110";
		Trees_din <= x"004134b5";
		wait for Clk_period;
		Addr <=  "0110100100111";
		Trees_din <= x"74000f04";
		wait for Clk_period;
		Addr <=  "0110100101000";
		Trees_din <= x"000b34b5";
		wait for Clk_period;
		Addr <=  "0110100101001";
		Trees_din <= x"ffd934b5";
		wait for Clk_period;
		Addr <=  "0110100101010";
		Trees_din <= x"82ff1a04";
		wait for Clk_period;
		Addr <=  "0110100101011";
		Trees_din <= x"fff934b5";
		wait for Clk_period;
		Addr <=  "0110100101100";
		Trees_din <= x"008934b5";
		wait for Clk_period;
		Addr <=  "0110100101101";
		Trees_din <= x"0700b158";
		wait for Clk_period;
		Addr <=  "0110100101110";
		Trees_din <= x"85003238";
		wait for Clk_period;
		Addr <=  "0110100101111";
		Trees_din <= x"2ffffe20";
		wait for Clk_period;
		Addr <=  "0110100110000";
		Trees_din <= x"7bff7f10";
		wait for Clk_period;
		Addr <=  "0110100110001";
		Trees_din <= x"a4ff8d08";
		wait for Clk_period;
		Addr <=  "0110100110010";
		Trees_din <= x"a5feb704";
		wait for Clk_period;
		Addr <=  "0110100110011";
		Trees_din <= x"ffd63609";
		wait for Clk_period;
		Addr <=  "0110100110100";
		Trees_din <= x"00233609";
		wait for Clk_period;
		Addr <=  "0110100110101";
		Trees_din <= x"d3ff5204";
		wait for Clk_period;
		Addr <=  "0110100110110";
		Trees_din <= x"ffe83609";
		wait for Clk_period;
		Addr <=  "0110100110111";
		Trees_din <= x"00433609";
		wait for Clk_period;
		Addr <=  "0110100111000";
		Trees_din <= x"b3ff8208";
		wait for Clk_period;
		Addr <=  "0110100111001";
		Trees_din <= x"81ff2b04";
		wait for Clk_period;
		Addr <=  "0110100111010";
		Trees_din <= x"00273609";
		wait for Clk_period;
		Addr <=  "0110100111011";
		Trees_din <= x"ffcf3609";
		wait for Clk_period;
		Addr <=  "0110100111100";
		Trees_din <= x"35ff4f04";
		wait for Clk_period;
		Addr <=  "0110100111101";
		Trees_din <= x"00513609";
		wait for Clk_period;
		Addr <=  "0110100111110";
		Trees_din <= x"ffba3609";
		wait for Clk_period;
		Addr <=  "0110100111111";
		Trees_din <= x"79feea0c";
		wait for Clk_period;
		Addr <=  "0110101000000";
		Trees_din <= x"befff504";
		wait for Clk_period;
		Addr <=  "0110101000001";
		Trees_din <= x"ffba3609";
		wait for Clk_period;
		Addr <=  "0110101000010";
		Trees_din <= x"6fff5904";
		wait for Clk_period;
		Addr <=  "0110101000011";
		Trees_din <= x"00803609";
		wait for Clk_period;
		Addr <=  "0110101000100";
		Trees_din <= x"fff33609";
		wait for Clk_period;
		Addr <=  "0110101000101";
		Trees_din <= x"bffffc08";
		wait for Clk_period;
		Addr <=  "0110101000110";
		Trees_din <= x"1dffa104";
		wait for Clk_period;
		Addr <=  "0110101000111";
		Trees_din <= x"ff793609";
		wait for Clk_period;
		Addr <=  "0110101001000";
		Trees_din <= x"00013609";
		wait for Clk_period;
		Addr <=  "0110101001001";
		Trees_din <= x"00203609";
		wait for Clk_period;
		Addr <=  "0110101001010";
		Trees_din <= x"26005b0c";
		wait for Clk_period;
		Addr <=  "0110101001011";
		Trees_din <= x"d5008908";
		wait for Clk_period;
		Addr <=  "0110101001100";
		Trees_din <= x"fe007f04";
		wait for Clk_period;
		Addr <=  "0110101001101";
		Trees_din <= x"ff6e3609";
		wait for Clk_period;
		Addr <=  "0110101001110";
		Trees_din <= x"00013609";
		wait for Clk_period;
		Addr <=  "0110101001111";
		Trees_din <= x"00163609";
		wait for Clk_period;
		Addr <=  "0110101010000";
		Trees_din <= x"30ff9a08";
		wait for Clk_period;
		Addr <=  "0110101010001";
		Trees_din <= x"3bff4a04";
		wait for Clk_period;
		Addr <=  "0110101010010";
		Trees_din <= x"ffe33609";
		wait for Clk_period;
		Addr <=  "0110101010011";
		Trees_din <= x"008a3609";
		wait for Clk_period;
		Addr <=  "0110101010100";
		Trees_din <= x"d4ff3708";
		wait for Clk_period;
		Addr <=  "0110101010101";
		Trees_din <= x"4cff3004";
		wait for Clk_period;
		Addr <=  "0110101010110";
		Trees_din <= x"ffb63609";
		wait for Clk_period;
		Addr <=  "0110101010111";
		Trees_din <= x"003d3609";
		wait for Clk_period;
		Addr <=  "0110101011000";
		Trees_din <= x"ff893609";
		wait for Clk_period;
		Addr <=  "0110101011001";
		Trees_din <= x"90fefc20";
		wait for Clk_period;
		Addr <=  "0110101011010";
		Trees_din <= x"1cff2e10";
		wait for Clk_period;
		Addr <=  "0110101011011";
		Trees_din <= x"33ff7a0c";
		wait for Clk_period;
		Addr <=  "0110101011100";
		Trees_din <= x"74000004";
		wait for Clk_period;
		Addr <=  "0110101011101";
		Trees_din <= x"007d3609";
		wait for Clk_period;
		Addr <=  "0110101011110";
		Trees_din <= x"69ff4704";
		wait for Clk_period;
		Addr <=  "0110101011111";
		Trees_din <= x"00393609";
		wait for Clk_period;
		Addr <=  "0110101100000";
		Trees_din <= x"ffa03609";
		wait for Clk_period;
		Addr <=  "0110101100001";
		Trees_din <= x"ffaa3609";
		wait for Clk_period;
		Addr <=  "0110101100010";
		Trees_din <= x"a4ffcc0c";
		wait for Clk_period;
		Addr <=  "0110101100011";
		Trees_din <= x"cf000604";
		wait for Clk_period;
		Addr <=  "0110101100100";
		Trees_din <= x"00143609";
		wait for Clk_period;
		Addr <=  "0110101100101";
		Trees_din <= x"a3ffb304";
		wait for Clk_period;
		Addr <=  "0110101100110";
		Trees_din <= x"00953609";
		wait for Clk_period;
		Addr <=  "0110101100111";
		Trees_din <= x"00133609";
		wait for Clk_period;
		Addr <=  "0110101101000";
		Trees_din <= x"ffe43609";
		wait for Clk_period;
		Addr <=  "0110101101001";
		Trees_din <= x"b9ff5320";
		wait for Clk_period;
		Addr <=  "0110101101010";
		Trees_din <= x"f5004410";
		wait for Clk_period;
		Addr <=  "0110101101011";
		Trees_din <= x"db00c808";
		wait for Clk_period;
		Addr <=  "0110101101100";
		Trees_din <= x"8b003704";
		wait for Clk_period;
		Addr <=  "0110101101101";
		Trees_din <= x"00383609";
		wait for Clk_period;
		Addr <=  "0110101101110";
		Trees_din <= x"ffda3609";
		wait for Clk_period;
		Addr <=  "0110101101111";
		Trees_din <= x"a3ff2304";
		wait for Clk_period;
		Addr <=  "0110101110000";
		Trees_din <= x"002f3609";
		wait for Clk_period;
		Addr <=  "0110101110001";
		Trees_din <= x"ffb73609";
		wait for Clk_period;
		Addr <=  "0110101110010";
		Trees_din <= x"7dff8b08";
		wait for Clk_period;
		Addr <=  "0110101110011";
		Trees_din <= x"d9ffa004";
		wait for Clk_period;
		Addr <=  "0110101110100";
		Trees_din <= x"ffbe3609";
		wait for Clk_period;
		Addr <=  "0110101110101";
		Trees_din <= x"00553609";
		wait for Clk_period;
		Addr <=  "0110101110110";
		Trees_din <= x"1dff6f04";
		wait for Clk_period;
		Addr <=  "0110101110111";
		Trees_din <= x"ff9b3609";
		wait for Clk_period;
		Addr <=  "0110101111000";
		Trees_din <= x"00273609";
		wait for Clk_period;
		Addr <=  "0110101111001";
		Trees_din <= x"d3ff6d10";
		wait for Clk_period;
		Addr <=  "0110101111010";
		Trees_din <= x"58ff5708";
		wait for Clk_period;
		Addr <=  "0110101111011";
		Trees_din <= x"c4feb804";
		wait for Clk_period;
		Addr <=  "0110101111100";
		Trees_din <= x"ffdf3609";
		wait for Clk_period;
		Addr <=  "0110101111101";
		Trees_din <= x"007b3609";
		wait for Clk_period;
		Addr <=  "0110101111110";
		Trees_din <= x"68fe8804";
		wait for Clk_period;
		Addr <=  "0110101111111";
		Trees_din <= x"00473609";
		wait for Clk_period;
		Addr <=  "0110110000000";
		Trees_din <= x"ffbe3609";
		wait for Clk_period;
		Addr <=  "0110110000001";
		Trees_din <= x"ffb83609";
		wait for Clk_period;
		Addr <=  "0110110000010";
		Trees_din <= x"0800c960";
		wait for Clk_period;
		Addr <=  "0110110000011";
		Trees_din <= x"6f003e40";
		wait for Clk_period;
		Addr <=  "0110110000100";
		Trees_din <= x"4cfeb420";
		wait for Clk_period;
		Addr <=  "0110110000101";
		Trees_din <= x"edffc810";
		wait for Clk_period;
		Addr <=  "0110110000110";
		Trees_din <= x"b2000308";
		wait for Clk_period;
		Addr <=  "0110110000111";
		Trees_din <= x"45ff3904";
		wait for Clk_period;
		Addr <=  "0110110001000";
		Trees_din <= x"ffaf375d";
		wait for Clk_period;
		Addr <=  "0110110001001";
		Trees_din <= x"0021375d";
		wait for Clk_period;
		Addr <=  "0110110001010";
		Trees_din <= x"e6ff7104";
		wait for Clk_period;
		Addr <=  "0110110001011";
		Trees_din <= x"ffa8375d";
		wait for Clk_period;
		Addr <=  "0110110001100";
		Trees_din <= x"003e375d";
		wait for Clk_period;
		Addr <=  "0110110001101";
		Trees_din <= x"0efdbd08";
		wait for Clk_period;
		Addr <=  "0110110001110";
		Trees_din <= x"91ff9e04";
		wait for Clk_period;
		Addr <=  "0110110001111";
		Trees_din <= x"0052375d";
		wait for Clk_period;
		Addr <=  "0110110010000";
		Trees_din <= x"ffbd375d";
		wait for Clk_period;
		Addr <=  "0110110010001";
		Trees_din <= x"e9ff9204";
		wait for Clk_period;
		Addr <=  "0110110010010";
		Trees_din <= x"ff71375d";
		wait for Clk_period;
		Addr <=  "0110110010011";
		Trees_din <= x"fff5375d";
		wait for Clk_period;
		Addr <=  "0110110010100";
		Trees_din <= x"60ff7c10";
		wait for Clk_period;
		Addr <=  "0110110010101";
		Trees_din <= x"e6002408";
		wait for Clk_period;
		Addr <=  "0110110010110";
		Trees_din <= x"78ffcb04";
		wait for Clk_period;
		Addr <=  "0110110010111";
		Trees_din <= x"0002375d";
		wait for Clk_period;
		Addr <=  "0110110011000";
		Trees_din <= x"ffbd375d";
		wait for Clk_period;
		Addr <=  "0110110011001";
		Trees_din <= x"33fe9904";
		wait for Clk_period;
		Addr <=  "0110110011010";
		Trees_din <= x"0046375d";
		wait for Clk_period;
		Addr <=  "0110110011011";
		Trees_din <= x"ff89375d";
		wait for Clk_period;
		Addr <=  "0110110011100";
		Trees_din <= x"6cff1008";
		wait for Clk_period;
		Addr <=  "0110110011101";
		Trees_din <= x"cdfff604";
		wait for Clk_period;
		Addr <=  "0110110011110";
		Trees_din <= x"0000375d";
		wait for Clk_period;
		Addr <=  "0110110011111";
		Trees_din <= x"ff91375d";
		wait for Clk_period;
		Addr <=  "0110110100000";
		Trees_din <= x"d3ff0b04";
		wait for Clk_period;
		Addr <=  "0110110100001";
		Trees_din <= x"0002375d";
		wait for Clk_period;
		Addr <=  "0110110100010";
		Trees_din <= x"0030375d";
		wait for Clk_period;
		Addr <=  "0110110100011";
		Trees_din <= x"f6fec108";
		wait for Clk_period;
		Addr <=  "0110110100100";
		Trees_din <= x"a9ffc404";
		wait for Clk_period;
		Addr <=  "0110110100101";
		Trees_din <= x"ffaf375d";
		wait for Clk_period;
		Addr <=  "0110110100110";
		Trees_din <= x"0031375d";
		wait for Clk_period;
		Addr <=  "0110110100111";
		Trees_din <= x"7aff5c0c";
		wait for Clk_period;
		Addr <=  "0110110101000";
		Trees_din <= x"90ff5808";
		wait for Clk_period;
		Addr <=  "0110110101001";
		Trees_din <= x"f202e204";
		wait for Clk_period;
		Addr <=  "0110110101010";
		Trees_din <= x"fffe375d";
		wait for Clk_period;
		Addr <=  "0110110101011";
		Trees_din <= x"0064375d";
		wait for Clk_period;
		Addr <=  "0110110101100";
		Trees_din <= x"ffad375d";
		wait for Clk_period;
		Addr <=  "0110110101101";
		Trees_din <= x"bfff6104";
		wait for Clk_period;
		Addr <=  "0110110101110";
		Trees_din <= x"fff7375d";
		wait for Clk_period;
		Addr <=  "0110110101111";
		Trees_din <= x"3f006104";
		wait for Clk_period;
		Addr <=  "0110110110000";
		Trees_din <= x"008a375d";
		wait for Clk_period;
		Addr <=  "0110110110001";
		Trees_din <= x"fff6375d";
		wait for Clk_period;
		Addr <=  "0110110110010";
		Trees_din <= x"5cffcd1c";
		wait for Clk_period;
		Addr <=  "0110110110011";
		Trees_din <= x"75fff910";
		wait for Clk_period;
		Addr <=  "0110110110100";
		Trees_din <= x"15ff9f08";
		wait for Clk_period;
		Addr <=  "0110110110101";
		Trees_din <= x"f0ff4b04";
		wait for Clk_period;
		Addr <=  "0110110110110";
		Trees_din <= x"007e375d";
		wait for Clk_period;
		Addr <=  "0110110110111";
		Trees_din <= x"fff7375d";
		wait for Clk_period;
		Addr <=  "0110110111000";
		Trees_din <= x"b3ff2204";
		wait for Clk_period;
		Addr <=  "0110110111001";
		Trees_din <= x"001a375d";
		wait for Clk_period;
		Addr <=  "0110110111010";
		Trees_din <= x"ff97375d";
		wait for Clk_period;
		Addr <=  "0110110111011";
		Trees_din <= x"0bfff604";
		wait for Clk_period;
		Addr <=  "0110110111100";
		Trees_din <= x"ff78375d";
		wait for Clk_period;
		Addr <=  "0110110111101";
		Trees_din <= x"a4ff7704";
		wait for Clk_period;
		Addr <=  "0110110111110";
		Trees_din <= x"ffa4375d";
		wait for Clk_period;
		Addr <=  "0110110111111";
		Trees_din <= x"0026375d";
		wait for Clk_period;
		Addr <=  "0110111000000";
		Trees_din <= x"8800c520";
		wait for Clk_period;
		Addr <=  "0110111000001";
		Trees_din <= x"48ff5310";
		wait for Clk_period;
		Addr <=  "0110111000010";
		Trees_din <= x"e2fe5508";
		wait for Clk_period;
		Addr <=  "0110111000011";
		Trees_din <= x"16fe9704";
		wait for Clk_period;
		Addr <=  "0110111000100";
		Trees_din <= x"fffa375d";
		wait for Clk_period;
		Addr <=  "0110111000101";
		Trees_din <= x"ff8d375d";
		wait for Clk_period;
		Addr <=  "0110111000110";
		Trees_din <= x"15ffb004";
		wait for Clk_period;
		Addr <=  "0110111000111";
		Trees_din <= x"ffe4375d";
		wait for Clk_period;
		Addr <=  "0110111001000";
		Trees_din <= x"0067375d";
		wait for Clk_period;
		Addr <=  "0110111001001";
		Trees_din <= x"62ff4908";
		wait for Clk_period;
		Addr <=  "0110111001010";
		Trees_din <= x"a0ff1d04";
		wait for Clk_period;
		Addr <=  "0110111001011";
		Trees_din <= x"007b375d";
		wait for Clk_period;
		Addr <=  "0110111001100";
		Trees_din <= x"000c375d";
		wait for Clk_period;
		Addr <=  "0110111001101";
		Trees_din <= x"b1ff0404";
		wait for Clk_period;
		Addr <=  "0110111001110";
		Trees_din <= x"0045375d";
		wait for Clk_period;
		Addr <=  "0110111001111";
		Trees_din <= x"ffd5375d";
		wait for Clk_period;
		Addr <=  "0110111010000";
		Trees_din <= x"91ff6b04";
		wait for Clk_period;
		Addr <=  "0110111010001";
		Trees_din <= x"0043375d";
		wait for Clk_period;
		Addr <=  "0110111010010";
		Trees_din <= x"ecffdd04";
		wait for Clk_period;
		Addr <=  "0110111010011";
		Trees_din <= x"001d375d";
		wait for Clk_period;
		Addr <=  "0110111010100";
		Trees_din <= x"1eff1304";
		wait for Clk_period;
		Addr <=  "0110111010101";
		Trees_din <= x"0006375d";
		wait for Clk_period;
		Addr <=  "0110111010110";
		Trees_din <= x"ff87375d";
		wait for Clk_period;
		Addr <=  "0110111010111";
		Trees_din <= x"d500a268";
		wait for Clk_period;
		Addr <=  "0110111011000";
		Trees_din <= x"7200472c";
		wait for Clk_period;
		Addr <=  "0110111011001";
		Trees_din <= x"65001a20";
		wait for Clk_period;
		Addr <=  "0110111011010";
		Trees_din <= x"b3ff9410";
		wait for Clk_period;
		Addr <=  "0110111011011";
		Trees_din <= x"1efef208";
		wait for Clk_period;
		Addr <=  "0110111011100";
		Trees_din <= x"60ffba04";
		wait for Clk_period;
		Addr <=  "0110111011101";
		Trees_din <= x"00073861";
		wait for Clk_period;
		Addr <=  "0110111011110";
		Trees_din <= x"00763861";
		wait for Clk_period;
		Addr <=  "0110111011111";
		Trees_din <= x"06ff7404";
		wait for Clk_period;
		Addr <=  "0110111100000";
		Trees_din <= x"00083861";
		wait for Clk_period;
		Addr <=  "0110111100001";
		Trees_din <= x"ffe13861";
		wait for Clk_period;
		Addr <=  "0110111100010";
		Trees_din <= x"55ffd708";
		wait for Clk_period;
		Addr <=  "0110111100011";
		Trees_din <= x"edffc504";
		wait for Clk_period;
		Addr <=  "0110111100100";
		Trees_din <= x"007d3861";
		wait for Clk_period;
		Addr <=  "0110111100101";
		Trees_din <= x"ffe13861";
		wait for Clk_period;
		Addr <=  "0110111100110";
		Trees_din <= x"b1ff2204";
		wait for Clk_period;
		Addr <=  "0110111100111";
		Trees_din <= x"ffdc3861";
		wait for Clk_period;
		Addr <=  "0110111101000";
		Trees_din <= x"003e3861";
		wait for Clk_period;
		Addr <=  "0110111101001";
		Trees_din <= x"6fffda08";
		wait for Clk_period;
		Addr <=  "0110111101010";
		Trees_din <= x"d3fea104";
		wait for Clk_period;
		Addr <=  "0110111101011";
		Trees_din <= x"ffec3861";
		wait for Clk_period;
		Addr <=  "0110111101100";
		Trees_din <= x"ff7a3861";
		wait for Clk_period;
		Addr <=  "0110111101101";
		Trees_din <= x"002b3861";
		wait for Clk_period;
		Addr <=  "0110111101110";
		Trees_din <= x"45fe7f20";
		wait for Clk_period;
		Addr <=  "0110111101111";
		Trees_din <= x"6e004910";
		wait for Clk_period;
		Addr <=  "0110111110000";
		Trees_din <= x"e1ffd908";
		wait for Clk_period;
		Addr <=  "0110111110001";
		Trees_din <= x"a1fe4204";
		wait for Clk_period;
		Addr <=  "0110111110010";
		Trees_din <= x"00043861";
		wait for Clk_period;
		Addr <=  "0110111110011";
		Trees_din <= x"ff733861";
		wait for Clk_period;
		Addr <=  "0110111110100";
		Trees_din <= x"2200c804";
		wait for Clk_period;
		Addr <=  "0110111110101";
		Trees_din <= x"ffbc3861";
		wait for Clk_period;
		Addr <=  "0110111110110";
		Trees_din <= x"004d3861";
		wait for Clk_period;
		Addr <=  "0110111110111";
		Trees_din <= x"05003208";
		wait for Clk_period;
		Addr <=  "0110111111000";
		Trees_din <= x"28ff2a04";
		wait for Clk_period;
		Addr <=  "0110111111001";
		Trees_din <= x"00003861";
		wait for Clk_period;
		Addr <=  "0110111111010";
		Trees_din <= x"ffa63861";
		wait for Clk_period;
		Addr <=  "0110111111011";
		Trees_din <= x"63ffc604";
		wait for Clk_period;
		Addr <=  "0110111111100";
		Trees_din <= x"005f3861";
		wait for Clk_period;
		Addr <=  "0110111111101";
		Trees_din <= x"ffd43861";
		wait for Clk_period;
		Addr <=  "0110111111110";
		Trees_din <= x"96fefd0c";
		wait for Clk_period;
		Addr <=  "0110111111111";
		Trees_din <= x"2bfeca04";
		wait for Clk_period;
		Addr <=  "0111000000000";
		Trees_din <= x"ffc23861";
		wait for Clk_period;
		Addr <=  "0111000000001";
		Trees_din <= x"16ff2204";
		wait for Clk_period;
		Addr <=  "0111000000010";
		Trees_din <= x"00763861";
		wait for Clk_period;
		Addr <=  "0111000000011";
		Trees_din <= x"00053861";
		wait for Clk_period;
		Addr <=  "0111000000100";
		Trees_din <= x"94ff9808";
		wait for Clk_period;
		Addr <=  "0111000000101";
		Trees_din <= x"11ff3b04";
		wait for Clk_period;
		Addr <=  "0111000000110";
		Trees_din <= x"004f3861";
		wait for Clk_period;
		Addr <=  "0111000000111";
		Trees_din <= x"00033861";
		wait for Clk_period;
		Addr <=  "0111000001000";
		Trees_din <= x"59ffae04";
		wait for Clk_period;
		Addr <=  "0111000001001";
		Trees_din <= x"00133861";
		wait for Clk_period;
		Addr <=  "0111000001010";
		Trees_din <= x"ffc73861";
		wait for Clk_period;
		Addr <=  "0111000001011";
		Trees_din <= x"af002118";
		wait for Clk_period;
		Addr <=  "0111000001100";
		Trees_din <= x"9bfeb404";
		wait for Clk_period;
		Addr <=  "0111000001101";
		Trees_din <= x"ffdc3861";
		wait for Clk_period;
		Addr <=  "0111000001110";
		Trees_din <= x"04009508";
		wait for Clk_period;
		Addr <=  "0111000001111";
		Trees_din <= x"e4feee04";
		wait for Clk_period;
		Addr <=  "0111000010000";
		Trees_din <= x"ffb03861";
		wait for Clk_period;
		Addr <=  "0111000010001";
		Trees_din <= x"005b3861";
		wait for Clk_period;
		Addr <=  "0111000010010";
		Trees_din <= x"e6ff4a04";
		wait for Clk_period;
		Addr <=  "0111000010011";
		Trees_din <= x"000f3861";
		wait for Clk_period;
		Addr <=  "0111000010100";
		Trees_din <= x"e0fec504";
		wait for Clk_period;
		Addr <=  "0111000010101";
		Trees_din <= x"002b3861";
		wait for Clk_period;
		Addr <=  "0111000010110";
		Trees_din <= x"00883861";
		wait for Clk_period;
		Addr <=  "0111000010111";
		Trees_din <= x"ffc53861";
		wait for Clk_period;
		Addr <=  "0111000011000";
		Trees_din <= x"25007850";
		wait for Clk_period;
		Addr <=  "0111000011001";
		Trees_din <= x"3cff7e38";
		wait for Clk_period;
		Addr <=  "0111000011010";
		Trees_din <= x"f1000c20";
		wait for Clk_period;
		Addr <=  "0111000011011";
		Trees_din <= x"2dff1510";
		wait for Clk_period;
		Addr <=  "0111000011100";
		Trees_din <= x"63ffec08";
		wait for Clk_period;
		Addr <=  "0111000011101";
		Trees_din <= x"40000404";
		wait for Clk_period;
		Addr <=  "0111000011110";
		Trees_din <= x"ffd739bd";
		wait for Clk_period;
		Addr <=  "0111000011111";
		Trees_din <= x"000239bd";
		wait for Clk_period;
		Addr <=  "0111000100000";
		Trees_din <= x"6affbe04";
		wait for Clk_period;
		Addr <=  "0111000100001";
		Trees_din <= x"fffe39bd";
		wait for Clk_period;
		Addr <=  "0111000100010";
		Trees_din <= x"004839bd";
		wait for Clk_period;
		Addr <=  "0111000100011";
		Trees_din <= x"01fec208";
		wait for Clk_period;
		Addr <=  "0111000100100";
		Trees_din <= x"00ff0504";
		wait for Clk_period;
		Addr <=  "0111000100101";
		Trees_din <= x"ffdf39bd";
		wait for Clk_period;
		Addr <=  "0111000100110";
		Trees_din <= x"003f39bd";
		wait for Clk_period;
		Addr <=  "0111000100111";
		Trees_din <= x"c1feb204";
		wait for Clk_period;
		Addr <=  "0111000101000";
		Trees_din <= x"ffc839bd";
		wait for Clk_period;
		Addr <=  "0111000101001";
		Trees_din <= x"001f39bd";
		wait for Clk_period;
		Addr <=  "0111000101010";
		Trees_din <= x"9bfeeb0c";
		wait for Clk_period;
		Addr <=  "0111000101011";
		Trees_din <= x"64fedf04";
		wait for Clk_period;
		Addr <=  "0111000101100";
		Trees_din <= x"ffa639bd";
		wait for Clk_period;
		Addr <=  "0111000101101";
		Trees_din <= x"b2ffde04";
		wait for Clk_period;
		Addr <=  "0111000101110";
		Trees_din <= x"006439bd";
		wait for Clk_period;
		Addr <=  "0111000101111";
		Trees_din <= x"ffd139bd";
		wait for Clk_period;
		Addr <=  "0111000110000";
		Trees_din <= x"c0ffbc08";
		wait for Clk_period;
		Addr <=  "0111000110001";
		Trees_din <= x"0800eb04";
		wait for Clk_period;
		Addr <=  "0111000110010";
		Trees_din <= x"ff8239bd";
		wait for Clk_period;
		Addr <=  "0111000110011";
		Trees_din <= x"000839bd";
		wait for Clk_period;
		Addr <=  "0111000110100";
		Trees_din <= x"002539bd";
		wait for Clk_period;
		Addr <=  "0111000110101";
		Trees_din <= x"b9fe9108";
		wait for Clk_period;
		Addr <=  "0111000110110";
		Trees_din <= x"49001504";
		wait for Clk_period;
		Addr <=  "0111000110111";
		Trees_din <= x"ffe739bd";
		wait for Clk_period;
		Addr <=  "0111000111000";
		Trees_din <= x"006739bd";
		wait for Clk_period;
		Addr <=  "0111000111001";
		Trees_din <= x"41ff6f08";
		wait for Clk_period;
		Addr <=  "0111000111010";
		Trees_din <= x"f6fea504";
		wait for Clk_period;
		Addr <=  "0111000111011";
		Trees_din <= x"000c39bd";
		wait for Clk_period;
		Addr <=  "0111000111100";
		Trees_din <= x"ff7839bd";
		wait for Clk_period;
		Addr <=  "0111000111101";
		Trees_din <= x"eeffdb04";
		wait for Clk_period;
		Addr <=  "0111000111110";
		Trees_din <= x"005f39bd";
		wait for Clk_period;
		Addr <=  "0111000111111";
		Trees_din <= x"ffc339bd";
		wait for Clk_period;
		Addr <=  "0111001000000";
		Trees_din <= x"5fff2b28";
		wait for Clk_period;
		Addr <=  "0111001000001";
		Trees_din <= x"5dff2108";
		wait for Clk_period;
		Addr <=  "0111001000010";
		Trees_din <= x"29ff5404";
		wait for Clk_period;
		Addr <=  "0111001000011";
		Trees_din <= x"000939bd";
		wait for Clk_period;
		Addr <=  "0111001000100";
		Trees_din <= x"ff8f39bd";
		wait for Clk_period;
		Addr <=  "0111001000101";
		Trees_din <= x"ccffad10";
		wait for Clk_period;
		Addr <=  "0111001000110";
		Trees_din <= x"bcfef708";
		wait for Clk_period;
		Addr <=  "0111001000111";
		Trees_din <= x"47ff9904";
		wait for Clk_period;
		Addr <=  "0111001001000";
		Trees_din <= x"ffe339bd";
		wait for Clk_period;
		Addr <=  "0111001001001";
		Trees_din <= x"006239bd";
		wait for Clk_period;
		Addr <=  "0111001001010";
		Trees_din <= x"a2000004";
		wait for Clk_period;
		Addr <=  "0111001001011";
		Trees_din <= x"ffb939bd";
		wait for Clk_period;
		Addr <=  "0111001001100";
		Trees_din <= x"004339bd";
		wait for Clk_period;
		Addr <=  "0111001001101";
		Trees_din <= x"2b00a508";
		wait for Clk_period;
		Addr <=  "0111001001110";
		Trees_din <= x"11ffb704";
		wait for Clk_period;
		Addr <=  "0111001001111";
		Trees_din <= x"006839bd";
		wait for Clk_period;
		Addr <=  "0111001010000";
		Trees_din <= x"ffea39bd";
		wait for Clk_period;
		Addr <=  "0111001010001";
		Trees_din <= x"c3004104";
		wait for Clk_period;
		Addr <=  "0111001010010";
		Trees_din <= x"ffa739bd";
		wait for Clk_period;
		Addr <=  "0111001010011";
		Trees_din <= x"003d39bd";
		wait for Clk_period;
		Addr <=  "0111001010100";
		Trees_din <= x"93ff6418";
		wait for Clk_period;
		Addr <=  "0111001010101";
		Trees_din <= x"b9ff5b0c";
		wait for Clk_period;
		Addr <=  "0111001010110";
		Trees_din <= x"47ff2804";
		wait for Clk_period;
		Addr <=  "0111001010111";
		Trees_din <= x"005439bd";
		wait for Clk_period;
		Addr <=  "0111001011000";
		Trees_din <= x"f1ff2404";
		wait for Clk_period;
		Addr <=  "0111001011001";
		Trees_din <= x"003c39bd";
		wait for Clk_period;
		Addr <=  "0111001011010";
		Trees_din <= x"ff9039bd";
		wait for Clk_period;
		Addr <=  "0111001011011";
		Trees_din <= x"d0006b08";
		wait for Clk_period;
		Addr <=  "0111001011100";
		Trees_din <= x"1cff3b04";
		wait for Clk_period;
		Addr <=  "0111001011101";
		Trees_din <= x"007b39bd";
		wait for Clk_period;
		Addr <=  "0111001011110";
		Trees_din <= x"001239bd";
		wait for Clk_period;
		Addr <=  "0111001011111";
		Trees_din <= x"ffc939bd";
		wait for Clk_period;
		Addr <=  "0111001100000";
		Trees_din <= x"0bffeb10";
		wait for Clk_period;
		Addr <=  "0111001100001";
		Trees_din <= x"5bff6708";
		wait for Clk_period;
		Addr <=  "0111001100010";
		Trees_din <= x"d3ff4204";
		wait for Clk_period;
		Addr <=  "0111001100011";
		Trees_din <= x"ffad39bd";
		wait for Clk_period;
		Addr <=  "0111001100100";
		Trees_din <= x"004d39bd";
		wait for Clk_period;
		Addr <=  "0111001100101";
		Trees_din <= x"24ffda04";
		wait for Clk_period;
		Addr <=  "0111001100110";
		Trees_din <= x"008039bd";
		wait for Clk_period;
		Addr <=  "0111001100111";
		Trees_din <= x"ffef39bd";
		wait for Clk_period;
		Addr <=  "0111001101000";
		Trees_din <= x"3bff8108";
		wait for Clk_period;
		Addr <=  "0111001101001";
		Trees_din <= x"0800b804";
		wait for Clk_period;
		Addr <=  "0111001101010";
		Trees_din <= x"ff8e39bd";
		wait for Clk_period;
		Addr <=  "0111001101011";
		Trees_din <= x"001a39bd";
		wait for Clk_period;
		Addr <=  "0111001101100";
		Trees_din <= x"fdff8104";
		wait for Clk_period;
		Addr <=  "0111001101101";
		Trees_din <= x"005939bd";
		wait for Clk_period;
		Addr <=  "0111001101110";
		Trees_din <= x"ffd739bd";
		wait for Clk_period;
		Addr <=  "0111001101111";
		Trees_din <= x"d2ff9a78";
		wait for Clk_period;
		Addr <=  "0111001110000";
		Trees_din <= x"aeff4340";
		wait for Clk_period;
		Addr <=  "0111001110001";
		Trees_din <= x"e6ff3420";
		wait for Clk_period;
		Addr <=  "0111001110010";
		Trees_din <= x"91ff7310";
		wait for Clk_period;
		Addr <=  "0111001110011";
		Trees_din <= x"96ff3c08";
		wait for Clk_period;
		Addr <=  "0111001110100";
		Trees_din <= x"2dfedc04";
		wait for Clk_period;
		Addr <=  "0111001110101";
		Trees_din <= x"fff73ac9";
		wait for Clk_period;
		Addr <=  "0111001110110";
		Trees_din <= x"00623ac9";
		wait for Clk_period;
		Addr <=  "0111001110111";
		Trees_din <= x"ceffbb04";
		wait for Clk_period;
		Addr <=  "0111001111000";
		Trees_din <= x"ffb43ac9";
		wait for Clk_period;
		Addr <=  "0111001111001";
		Trees_din <= x"000e3ac9";
		wait for Clk_period;
		Addr <=  "0111001111010";
		Trees_din <= x"37fed108";
		wait for Clk_period;
		Addr <=  "0111001111011";
		Trees_din <= x"b9fee904";
		wait for Clk_period;
		Addr <=  "0111001111100";
		Trees_din <= x"ffd83ac9";
		wait for Clk_period;
		Addr <=  "0111001111101";
		Trees_din <= x"00483ac9";
		wait for Clk_period;
		Addr <=  "0111001111110";
		Trees_din <= x"f800c104";
		wait for Clk_period;
		Addr <=  "0111001111111";
		Trees_din <= x"ff893ac9";
		wait for Clk_period;
		Addr <=  "0111010000000";
		Trees_din <= x"000e3ac9";
		wait for Clk_period;
		Addr <=  "0111010000001";
		Trees_din <= x"72006910";
		wait for Clk_period;
		Addr <=  "0111010000010";
		Trees_din <= x"7efdfc08";
		wait for Clk_period;
		Addr <=  "0111010000011";
		Trees_din <= x"79ff5e04";
		wait for Clk_period;
		Addr <=  "0111010000100";
		Trees_din <= x"006b3ac9";
		wait for Clk_period;
		Addr <=  "0111010000101";
		Trees_din <= x"fff03ac9";
		wait for Clk_period;
		Addr <=  "0111010000110";
		Trees_din <= x"65001a04";
		wait for Clk_period;
		Addr <=  "0111010000111";
		Trees_din <= x"00023ac9";
		wait for Clk_period;
		Addr <=  "0111010001000";
		Trees_din <= x"ffab3ac9";
		wait for Clk_period;
		Addr <=  "0111010001001";
		Trees_din <= x"61ff6c08";
		wait for Clk_period;
		Addr <=  "0111010001010";
		Trees_din <= x"88ffd304";
		wait for Clk_period;
		Addr <=  "0111010001011";
		Trees_din <= x"ff983ac9";
		wait for Clk_period;
		Addr <=  "0111010001100";
		Trees_din <= x"00163ac9";
		wait for Clk_period;
		Addr <=  "0111010001101";
		Trees_din <= x"46fec704";
		wait for Clk_period;
		Addr <=  "0111010001110";
		Trees_din <= x"00043ac9";
		wait for Clk_period;
		Addr <=  "0111010001111";
		Trees_din <= x"00603ac9";
		wait for Clk_period;
		Addr <=  "0111010010000";
		Trees_din <= x"03ffb11c";
		wait for Clk_period;
		Addr <=  "0111010010001";
		Trees_din <= x"adffb50c";
		wait for Clk_period;
		Addr <=  "0111010010010";
		Trees_din <= x"f7fe8204";
		wait for Clk_period;
		Addr <=  "0111010010011";
		Trees_din <= x"00513ac9";
		wait for Clk_period;
		Addr <=  "0111010010100";
		Trees_din <= x"4900ab04";
		wait for Clk_period;
		Addr <=  "0111010010101";
		Trees_din <= x"ff983ac9";
		wait for Clk_period;
		Addr <=  "0111010010110";
		Trees_din <= x"00403ac9";
		wait for Clk_period;
		Addr <=  "0111010010111";
		Trees_din <= x"46ff0b08";
		wait for Clk_period;
		Addr <=  "0111010011000";
		Trees_din <= x"19ff6e04";
		wait for Clk_period;
		Addr <=  "0111010011001";
		Trees_din <= x"004d3ac9";
		wait for Clk_period;
		Addr <=  "0111010011010";
		Trees_din <= x"ffbb3ac9";
		wait for Clk_period;
		Addr <=  "0111010011011";
		Trees_din <= x"ebff1404";
		wait for Clk_period;
		Addr <=  "0111010011100";
		Trees_din <= x"ff953ac9";
		wait for Clk_period;
		Addr <=  "0111010011101";
		Trees_din <= x"fff63ac9";
		wait for Clk_period;
		Addr <=  "0111010011110";
		Trees_din <= x"0cfde20c";
		wait for Clk_period;
		Addr <=  "0111010011111";
		Trees_din <= x"47ffbb04";
		wait for Clk_period;
		Addr <=  "0111010100000";
		Trees_din <= x"ffad3ac9";
		wait for Clk_period;
		Addr <=  "0111010100001";
		Trees_din <= x"7eff0c04";
		wait for Clk_period;
		Addr <=  "0111010100010";
		Trees_din <= x"00813ac9";
		wait for Clk_period;
		Addr <=  "0111010100011";
		Trees_din <= x"ffe13ac9";
		wait for Clk_period;
		Addr <=  "0111010100100";
		Trees_din <= x"34fff508";
		wait for Clk_period;
		Addr <=  "0111010100101";
		Trees_din <= x"d600e604";
		wait for Clk_period;
		Addr <=  "0111010100110";
		Trees_din <= x"ffa73ac9";
		wait for Clk_period;
		Addr <=  "0111010100111";
		Trees_din <= x"00403ac9";
		wait for Clk_period;
		Addr <=  "0111010101000";
		Trees_din <= x"40fff704";
		wait for Clk_period;
		Addr <=  "0111010101001";
		Trees_din <= x"ffda3ac9";
		wait for Clk_period;
		Addr <=  "0111010101010";
		Trees_din <= x"00273ac9";
		wait for Clk_period;
		Addr <=  "0111010101011";
		Trees_din <= x"fdff4204";
		wait for Clk_period;
		Addr <=  "0111010101100";
		Trees_din <= x"ffdc3ac9";
		wait for Clk_period;
		Addr <=  "0111010101101";
		Trees_din <= x"b4ff5608";
		wait for Clk_period;
		Addr <=  "0111010101110";
		Trees_din <= x"36ff9504";
		wait for Clk_period;
		Addr <=  "0111010101111";
		Trees_din <= x"00893ac9";
		wait for Clk_period;
		Addr <=  "0111010110000";
		Trees_din <= x"00233ac9";
		wait for Clk_period;
		Addr <=  "0111010110001";
		Trees_din <= x"00093ac9";
		wait for Clk_period;
		Addr <=  "0111010110010";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  2
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"57002150";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"35fff930";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"9f004b20";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"f7012410";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"f6fe0c08";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"ceff7004";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"015e00dd";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"ffac00dd";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"b9002804";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"ff6d00dd";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"012800dd";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"b3fea108";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"2bff6704";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"003700dd";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"036600dd";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"e5fde304";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"01ef00dd";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"ff9100dd";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"dafff308";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"02feb504";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"00a600dd";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"036400dd";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"01fe6404";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"003700dd";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"ff9000dd";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"49ff7808";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"08008204";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"038700dd";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"ffa400dd";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"c4ff2f0c";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"2bffeb08";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"f7007f04";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"ffe800dd";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"030400dd";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"ff7c00dd";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"fb001908";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"41ff6904";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"ff6100dd";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"003700dd";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"010200dd";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"feff6608";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"07ffc004";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"003700dd";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"ff7900dd";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"56ff3a0c";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"65ff3f04";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"022f00dd";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"02fe4704";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"003700dd";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"ff8100dd";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"07ffd304";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"003700dd";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"8ffea704";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"003700dd";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"03e700dd";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"57000660";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"35ffc434";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"9f003f20";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"f7012410";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"f6fe0c08";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"f2024204";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"014b01e1";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"ff6a01e1";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"7b002d04";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"ff6f01e1";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"001201e1";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"88fffd08";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"b3ff4104";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"01cb01e1";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"ff9e01e1";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"d0ffda04";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"00d301e1";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"ff6a01e1";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"8800250c";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"ddff5408";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"f2026104";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"022401e1";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"000801e1";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"ff9e01e1";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"58fe9f04";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"003c01e1";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"ff8201e1";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"f700a118";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"7cff7010";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"f1fff908";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"6cfef004";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"00c801e1";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"ff6901e1";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"24ff6204";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"ff9f01e1";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"020d01e1";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"86ffe404";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"ff5d01e1";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"003b01e1";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"2a00ae10";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"39ffa008";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"96ff3104";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"004b01e1";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"023601e1";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"5a00a304";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"ff7901e1";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"00f201e1";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"ff7b01e1";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"beff2a0c";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"d8ffdf04";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"002101e1";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"b2ffe604";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"02bf01e1";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"00c301e1";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"8ffead04";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"ff6d01e1";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"feff6804";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"ff7801e1";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"83ff5708";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"a2ffa004";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"ff9d01e1";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"01dc01e1";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"0fff4004";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"00c201e1";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"ff7901e1";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"57ffc664";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"35ffc434";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"9f003f20";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"f7010f10";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"b9002808";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"d4ff9a04";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"ff6b031d";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"ffb2031d";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"d0002c04";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"ff8b031d";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"027c031d";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"e3fe4508";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"22004e04";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"0189031d";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"ffa1031d";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"1afe1d04";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"00f7031d";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"ff68031d";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"5bff6208";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"3cff0d04";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"0194031d";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"0018031d";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"c7ff6808";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"37001d04";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"ff77031d";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"0031031d";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"0100031d";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"b3fea114";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"a0ff2408";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"ddffb304";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"ff79031d";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"011d031d";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"78fed304";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"ffa2031d";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"33fef404";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"0009031d";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"01a8031d";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"cafeb60c";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"dcfedb04";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"0137031d";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"b6ffc904";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"ff5d031d";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"0043031d";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"abfffd08";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"a6ff6f04";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"0133031d";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"ff8e031d";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"47ff6d04";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"00ae031d";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"ff6e031d";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"beff3218";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"20ff0b04";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"ff9b031d";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"61feda0c";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"8dfe9a04";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"007f031d";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"73005904";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"021d031d";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"008f031d";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"45feb804";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"012c031d";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"ff8c031d";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"49ffb010";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"12ff2e04";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"ff75031d";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"71ff5f04";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"ff8e031d";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"d2fed204";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"0024031d";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"0201031d";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"6bfe3108";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"24ffc904";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"ffa0031d";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"013a031d";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"5dff0304";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"00ce031d";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"78ff0804";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"005d031d";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"ff6a031d";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"57ffc65c";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"35ffc434";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"9f003f20";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"7b002d10";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"a1ff2808";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"a6fe9d04";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"ffe70449";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"ff5f0449";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"f6fe5504";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"00730449";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"ff990449";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"3cff4208";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"5a00f304";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"ff660449";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"00be0449";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"49ffd104";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"01e30449";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"ff870449";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"c7ff680c";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"0bffa804";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"ff7f0449";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"19ff7304";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"ffd70449";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"01120449";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"56ff1b04";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"00630449";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"016a0449";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"b3feea14";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"2a009a0c";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"c2ffc808";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"2b003f04";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"010a0449";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"ff9c0449";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"ff8d0449";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"27fff104";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"ff7c0449";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"003c0449";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"0bfffd08";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"1cfe9a04";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"002c0449";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"ff620449";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"b6ff8008";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"b6ff4a04";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"ff950449";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"014c0449";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"ff7e0449";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"f6fee024";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"53ff7508";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"8effaa04";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"00d80449";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"ff700449";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"d2feb00c";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"e0ff2808";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"88002004";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"011c0449";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"ffa20449";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"ff790449";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"15ffb008";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"38ffaf04";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"01a90449";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"00430449";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"1b001104";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"ff890449";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"00cf0449";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"57002108";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"edff3504";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"00400449";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"ff650449";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"8bffea08";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"c7ff6704";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"00140449";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"01240449";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"faffc604";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"ff850449";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"00180449";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"f2026164";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"f6fe682c";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"c7feff0c";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"33ffdc08";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"daff5604";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"004e056d";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"ff67056d";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"00fa056d";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"93ff7910";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"ecffe008";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"db007e04";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"ff77056d";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"0029056d";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"7bff2504";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"0133056d";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"ff97056d";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"24ffd308";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"1bffb404";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"ff8e056d";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"00ea056d";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"8cffa304";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"031b056d";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"0115056d";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"f7009b1c";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"41ff390c";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"fdfe0504";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"0159056d";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"57001204";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"ff7d056d";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"005b056d";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"cbff7508";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"96001d04";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"002b056d";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"01fe056d";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"fcffd004";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"ffaa056d";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"00ab056d";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"2a007e0c";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"1dfeaa04";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"ff8a056d";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"f0ff6b04";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"011f056d";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"004e056d";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"59004e08";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"42feaa04";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"0020056d";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"ff65056d";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"00ff3404";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"00b8056d";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"0001056d";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"6dff8f08";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"d8008204";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"ff79056d";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"01ca056d";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"b3fe6110";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"b4ff2b08";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"0a015804";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"ff6e056d";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"0029056d";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"c8ffc704";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"0158056d";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"0008056d";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"f7014e10";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"7afed908";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"26fff804";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"014e056d";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"ff7c056d";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"c1fe0c04";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"002c056d";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"ff60056d";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"35ffa904";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"ffa8056d";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"00e7056d";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"f2026154";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"f6fe681c";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"24ff7208";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"c3005c04";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"ff730689";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"00140689";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"8dfe7204";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"ff7d0689";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"18ffd308";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"dcff9104";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"ffdf0689";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"01340689";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"d2febc04";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"ff7c0689";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"009b0689";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"e3fe541c";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"2a004f0c";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"23000408";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"afff1d04";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"01640689";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"00690689";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"ff740689";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"35000b08";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"5dff3c04";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"008c0689";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"ff670689";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"d0006304";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"ffac0689";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"01010689";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"49ffa510";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"8dff2608";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"43ffdb04";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"ff980689";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"007f0689";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"3bff6d04";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"00c30689";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"ff920689";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"5aff2004";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"01770689";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"57001204";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"ff840689";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"00500689";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"14ffac30";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"9fffb918";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"fdfe2f08";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"91ffa804";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"00d00689";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"ffac0689";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"7afe8d08";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"d1ff2904";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"ffa30689";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"00d40689";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"4ffe5e04";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"00010689";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"ff600689";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"55ff8708";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"47ffb404";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"01390689";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"ffa60689";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"d8008f08";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"d9ff5404";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"00310689";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"ff640689";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"5a008d04";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"ff990689";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"012d0689";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"6bff2008";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"31ff0f04";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"00460689";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"ff770689";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"017c0689";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"a1ff2830";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"7b002d24";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"9f004b1c";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"57ffc610";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"a6feb208";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"edff6e04";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"00be07cd";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"ff7807cd";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"8dff5404";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"ff6607cd";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"ffe107cd";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"24ffd304";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"ff7c07cd";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"6bfea604";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"00ee07cd";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"ffa007cd";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"07006f04";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"fffe07cd";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"00ca07cd";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"b9ff0e04";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"ff7e07cd";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"fdff9704";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"01af07cd";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"000707cd";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"16ff0c38";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"d3fe9518";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"47003010";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"96ff3f08";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"0dff8f04";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"ff8307cd";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"fff907cd";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"c1fee904";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"011c07cd";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"ff8a07cd";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"c4fe8d04";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"007a07cd";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"ff6e07cd";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"f6fe4010";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"19ffb308";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"a1fff104";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"ff8607cd";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"007a07cd";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"29ff4404";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"014207cd";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"004007cd";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"35ffd908";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"8cfe8a04";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"009307cd";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"ff6807cd";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"c4ff5504";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"00aa07cd";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"ff8007cd";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"f6fea61c";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"61ff7210";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"14ff3008";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"57ff8a04";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"ff9507cd";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"00b207cd";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"b5fe9204";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"ffc607cd";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"017b07cd";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"21ff8908";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"25002b04";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"ff9a07cd";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"010107cd";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"ff7507cd";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"35ff5b10";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"39fff908";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"06008704";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"ff8f07cd";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"00f307cd";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"0fff2804";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"013b07cd";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"ffd907cd";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"2a00ae08";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"68fea604";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"012807cd";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"004807cd";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"1eff1904";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"001007cd";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"ff7507cd";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"f202666c";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"41ff2b34";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"9fffc418";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"2c008d10";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"35ffcc08";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"96006104";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"ff8b0911";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"00c80911";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"c8ffc804";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"008d0911";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"ffa70911";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"67ff4404";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"ffc50911";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"01520911";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"beff6810";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"18ffb308";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"01feec04";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"002b0911";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"012a0911";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"e6ff9704";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"00280911";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"ff940911";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"6dff9a04";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"01070911";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"6fff4d04";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"00320911";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"ff690911";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"47003220";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"3afed510";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"c1ff0a08";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"8dfe4704";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"ffaf0911";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"017a0911";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"fcff0b04";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"00370911";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"ff8b0911";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"18ffa308";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"38ff9104";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"00c70911";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"fff00911";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"5aff9a04";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"00fb0911";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"ffc50911";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"27004b0c";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"35001608";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"54ff5504";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"00000911";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"ff640911";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"004a0911";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"16ff4a04";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"ff920911";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"05000904";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"01740911";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"00300911";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"14ffac2c";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"e3fdfa0c";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"f5005808";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"2500cd04";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"ff830911";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"00360911";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"00d10911";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"7afed910";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"73ff8308";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"10ff6504";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"01680911";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"001d0911";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"c9004204";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"ff760911";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"00090911";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"f1002208";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"35005d04";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"ff610911";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"00540911";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"4dfec104";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"ff7a0911";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"00650911";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"e5feae08";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"dbffc304";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"01cc0911";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"ffeb0911";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"ff7e0911";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"f2026670";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"6cff643c";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"18ffbb1c";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"f0ff930c";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"2a00ae08";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"12005704";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"00bc0a55";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"ff840a55";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"ff7a0a55";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"a4ffa608";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"1301d904";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"ff750a55";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"00810a55";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"1eff9404";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"ff8f0a55";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"00b00a55";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"a3ffcf10";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"02ff6908";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"83feaf04";
		wait for Clk_period;
		Addr <=  "0001001010111";
		Trees_din <= x"00350a55";
		wait for Clk_period;
		Addr <=  "0001001011000";
		Trees_din <= x"ff780a55";
		wait for Clk_period;
		Addr <=  "0001001011001";
		Trees_din <= x"e3fed604";
		wait for Clk_period;
		Addr <=  "0001001011010";
		Trees_din <= x"00a50a55";
		wait for Clk_period;
		Addr <=  "0001001011011";
		Trees_din <= x"ff7e0a55";
		wait for Clk_period;
		Addr <=  "0001001011100";
		Trees_din <= x"16ff0c08";
		wait for Clk_period;
		Addr <=  "0001001011101";
		Trees_din <= x"2a001104";
		wait for Clk_period;
		Addr <=  "0001001011110";
		Trees_din <= x"ff7c0a55";
		wait for Clk_period;
		Addr <=  "0001001011111";
		Trees_din <= x"fff60a55";
		wait for Clk_period;
		Addr <=  "0001001100000";
		Trees_din <= x"81ff5d04";
		wait for Clk_period;
		Addr <=  "0001001100001";
		Trees_din <= x"018a0a55";
		wait for Clk_period;
		Addr <=  "0001001100010";
		Trees_din <= x"001b0a55";
		wait for Clk_period;
		Addr <=  "0001001100011";
		Trees_din <= x"64ff251c";
		wait for Clk_period;
		Addr <=  "0001001100100";
		Trees_din <= x"b3fed20c";
		wait for Clk_period;
		Addr <=  "0001001100101";
		Trees_din <= x"9dffd308";
		wait for Clk_period;
		Addr <=  "0001001100110";
		Trees_din <= x"7efe5f04";
		wait for Clk_period;
		Addr <=  "0001001100111";
		Trees_din <= x"ff7f0a55";
		wait for Clk_period;
		Addr <=  "0001001101000";
		Trees_din <= x"00ac0a55";
		wait for Clk_period;
		Addr <=  "0001001101001";
		Trees_din <= x"ff7a0a55";
		wait for Clk_period;
		Addr <=  "0001001101010";
		Trees_din <= x"5ffe8f08";
		wait for Clk_period;
		Addr <=  "0001001101011";
		Trees_din <= x"b9ff6204";
		wait for Clk_period;
		Addr <=  "0001001101100";
		Trees_din <= x"ffdc0a55";
		wait for Clk_period;
		Addr <=  "0001001101101";
		Trees_din <= x"01600a55";
		wait for Clk_period;
		Addr <=  "0001001101110";
		Trees_din <= x"c2fe9004";
		wait for Clk_period;
		Addr <=  "0001001101111";
		Trees_din <= x"00480a55";
		wait for Clk_period;
		Addr <=  "0001001110000";
		Trees_din <= x"ff830a55";
		wait for Clk_period;
		Addr <=  "0001001110001";
		Trees_din <= x"57000610";
		wait for Clk_period;
		Addr <=  "0001001110010";
		Trees_din <= x"f6fe4b08";
		wait for Clk_period;
		Addr <=  "0001001110011";
		Trees_din <= x"cafdee04";
		wait for Clk_period;
		Addr <=  "0001001110100";
		Trees_din <= x"00d10a55";
		wait for Clk_period;
		Addr <=  "0001001110101";
		Trees_din <= x"ffa50a55";
		wait for Clk_period;
		Addr <=  "0001001110110";
		Trees_din <= x"4ffe7004";
		wait for Clk_period;
		Addr <=  "0001001110111";
		Trees_din <= x"002e0a55";
		wait for Clk_period;
		Addr <=  "0001001111000";
		Trees_din <= x"ff620a55";
		wait for Clk_period;
		Addr <=  "0001001111001";
		Trees_din <= x"60ff5d04";
		wait for Clk_period;
		Addr <=  "0001001111010";
		Trees_din <= x"00d70a55";
		wait for Clk_period;
		Addr <=  "0001001111011";
		Trees_din <= x"ffd00a55";
		wait for Clk_period;
		Addr <=  "0001001111100";
		Trees_din <= x"a1ff6014";
		wait for Clk_period;
		Addr <=  "0001001111101";
		Trees_din <= x"68fdd504";
		wait for Clk_period;
		Addr <=  "0001001111110";
		Trees_din <= x"002c0a55";
		wait for Clk_period;
		Addr <=  "0001001111111";
		Trees_din <= x"7b005e0c";
		wait for Clk_period;
		Addr <=  "0001010000000";
		Trees_din <= x"fa005208";
		wait for Clk_period;
		Addr <=  "0001010000001";
		Trees_din <= x"9afe7504";
		wait for Clk_period;
		Addr <=  "0001010000010";
		Trees_din <= x"fff90a55";
		wait for Clk_period;
		Addr <=  "0001010000011";
		Trees_din <= x"ff630a55";
		wait for Clk_period;
		Addr <=  "0001010000100";
		Trees_din <= x"fffc0a55";
		wait for Clk_period;
		Addr <=  "0001010000101";
		Trees_din <= x"002f0a55";
		wait for Clk_period;
		Addr <=  "0001010000110";
		Trees_din <= x"bd00b71c";
		wait for Clk_period;
		Addr <=  "0001010000111";
		Trees_din <= x"f4ff2610";
		wait for Clk_period;
		Addr <=  "0001010001000";
		Trees_din <= x"35ffe008";
		wait for Clk_period;
		Addr <=  "0001010001001";
		Trees_din <= x"3bfe6b04";
		wait for Clk_period;
		Addr <=  "0001010001010";
		Trees_din <= x"002b0a55";
		wait for Clk_period;
		Addr <=  "0001010001011";
		Trees_din <= x"ff660a55";
		wait for Clk_period;
		Addr <=  "0001010001100";
		Trees_din <= x"75004904";
		wait for Clk_period;
		Addr <=  "0001010001101";
		Trees_din <= x"ffad0a55";
		wait for Clk_period;
		Addr <=  "0001010001110";
		Trees_din <= x"00a30a55";
		wait for Clk_period;
		Addr <=  "0001010001111";
		Trees_din <= x"ac003e04";
		wait for Clk_period;
		Addr <=  "0001010010000";
		Trees_din <= x"ff7b0a55";
		wait for Clk_period;
		Addr <=  "0001010010001";
		Trees_din <= x"22005c04";
		wait for Clk_period;
		Addr <=  "0001010010010";
		Trees_din <= x"00fa0a55";
		wait for Clk_period;
		Addr <=  "0001010010011";
		Trees_din <= x"ff990a55";
		wait for Clk_period;
		Addr <=  "0001010010100";
		Trees_din <= x"01060a55";
		wait for Clk_period;
		Addr <=  "0001010010101";
		Trees_din <= x"f2026860";
		wait for Clk_period;
		Addr <=  "0001010010110";
		Trees_din <= x"4700443c";
		wait for Clk_period;
		Addr <=  "0001010010111";
		Trees_din <= x"3afeda1c";
		wait for Clk_period;
		Addr <=  "0001010011000";
		Trees_din <= x"c1fed710";
		wait for Clk_period;
		Addr <=  "0001010011001";
		Trees_din <= x"91ffde08";
		wait for Clk_period;
		Addr <=  "0001010011010";
		Trees_din <= x"e5ff0b04";
		wait for Clk_period;
		Addr <=  "0001010011011";
		Trees_din <= x"01160b89";
		wait for Clk_period;
		Addr <=  "0001010011100";
		Trees_din <= x"fff70b89";
		wait for Clk_period;
		Addr <=  "0001010011101";
		Trees_din <= x"2dfed404";
		wait for Clk_period;
		Addr <=  "0001010011110";
		Trees_din <= x"008d0b89";
		wait for Clk_period;
		Addr <=  "0001010011111";
		Trees_din <= x"ff880b89";
		wait for Clk_period;
		Addr <=  "0001010100000";
		Trees_din <= x"7bff5104";
		wait for Clk_period;
		Addr <=  "0001010100001";
		Trees_din <= x"ff750b89";
		wait for Clk_period;
		Addr <=  "0001010100010";
		Trees_din <= x"f6fef104";
		wait for Clk_period;
		Addr <=  "0001010100011";
		Trees_din <= x"00bb0b89";
		wait for Clk_period;
		Addr <=  "0001010100100";
		Trees_din <= x"ff8c0b89";
		wait for Clk_period;
		Addr <=  "0001010100101";
		Trees_din <= x"09fec010";
		wait for Clk_period;
		Addr <=  "0001010100110";
		Trees_din <= x"42ff6c08";
		wait for Clk_period;
		Addr <=  "0001010100111";
		Trees_din <= x"9fffb004";
		wait for Clk_period;
		Addr <=  "0001010101000";
		Trees_din <= x"ffac0b89";
		wait for Clk_period;
		Addr <=  "0001010101001";
		Trees_din <= x"00880b89";
		wait for Clk_period;
		Addr <=  "0001010101010";
		Trees_din <= x"23ffbd04";
		wait for Clk_period;
		Addr <=  "0001010101011";
		Trees_din <= x"011c0b89";
		wait for Clk_period;
		Addr <=  "0001010101100";
		Trees_din <= x"ffcf0b89";
		wait for Clk_period;
		Addr <=  "0001010101101";
		Trees_din <= x"61ff8108";
		wait for Clk_period;
		Addr <=  "0001010101110";
		Trees_din <= x"41ff2e04";
		wait for Clk_period;
		Addr <=  "0001010101111";
		Trees_din <= x"ffc80b89";
		wait for Clk_period;
		Addr <=  "0001010110000";
		Trees_din <= x"005b0b89";
		wait for Clk_period;
		Addr <=  "0001010110001";
		Trees_din <= x"f700c704";
		wait for Clk_period;
		Addr <=  "0001010110010";
		Trees_din <= x"ff880b89";
		wait for Clk_period;
		Addr <=  "0001010110011";
		Trees_din <= x"005b0b89";
		wait for Clk_period;
		Addr <=  "0001010110100";
		Trees_din <= x"f1002714";
		wait for Clk_period;
		Addr <=  "0001010110101";
		Trees_din <= x"fcffee0c";
		wait for Clk_period;
		Addr <=  "0001010110110";
		Trees_din <= x"a0fff808";
		wait for Clk_period;
		Addr <=  "0001010110111";
		Trees_din <= x"f7012404";
		wait for Clk_period;
		Addr <=  "0001010111000";
		Trees_din <= x"ff640b89";
		wait for Clk_period;
		Addr <=  "0001010111001";
		Trees_din <= x"00050b89";
		wait for Clk_period;
		Addr <=  "0001010111010";
		Trees_din <= x"003c0b89";
		wait for Clk_period;
		Addr <=  "0001010111011";
		Trees_din <= x"06001f04";
		wait for Clk_period;
		Addr <=  "0001010111100";
		Trees_din <= x"ff9d0b89";
		wait for Clk_period;
		Addr <=  "0001010111101";
		Trees_din <= x"00f70b89";
		wait for Clk_period;
		Addr <=  "0001010111110";
		Trees_din <= x"16ff2904";
		wait for Clk_period;
		Addr <=  "0001010111111";
		Trees_din <= x"ff880b89";
		wait for Clk_period;
		Addr <=  "0001011000000";
		Trees_din <= x"25002f08";
		wait for Clk_period;
		Addr <=  "0001011000001";
		Trees_din <= x"54002a04";
		wait for Clk_period;
		Addr <=  "0001011000010";
		Trees_din <= x"002f0b89";
		wait for Clk_period;
		Addr <=  "0001011000011";
		Trees_din <= x"00fa0b89";
		wait for Clk_period;
		Addr <=  "0001011000100";
		Trees_din <= x"ffda0b89";
		wait for Clk_period;
		Addr <=  "0001011000101";
		Trees_din <= x"a1ff6014";
		wait for Clk_period;
		Addr <=  "0001011000110";
		Trees_din <= x"9a00930c";
		wait for Clk_period;
		Addr <=  "0001011000111";
		Trees_din <= x"fa005208";
		wait for Clk_period;
		Addr <=  "0001011001000";
		Trees_din <= x"77007504";
		wait for Clk_period;
		Addr <=  "0001011001001";
		Trees_din <= x"ff640b89";
		wait for Clk_period;
		Addr <=  "0001011001010";
		Trees_din <= x"fff60b89";
		wait for Clk_period;
		Addr <=  "0001011001011";
		Trees_din <= x"00020b89";
		wait for Clk_period;
		Addr <=  "0001011001100";
		Trees_din <= x"09ff1d04";
		wait for Clk_period;
		Addr <=  "0001011001101";
		Trees_din <= x"00c10b89";
		wait for Clk_period;
		Addr <=  "0001011001110";
		Trees_din <= x"ffa40b89";
		wait for Clk_period;
		Addr <=  "0001011001111";
		Trees_din <= x"95ffd218";
		wait for Clk_period;
		Addr <=  "0001011010000";
		Trees_din <= x"f4ff610c";
		wait for Clk_period;
		Addr <=  "0001011010001";
		Trees_din <= x"b3fe3c04";
		wait for Clk_period;
		Addr <=  "0001011010010";
		Trees_din <= x"007f0b89";
		wait for Clk_period;
		Addr <=  "0001011010011";
		Trees_din <= x"36004804";
		wait for Clk_period;
		Addr <=  "0001011010100";
		Trees_din <= x"ff680b89";
		wait for Clk_period;
		Addr <=  "0001011010101";
		Trees_din <= x"00040b89";
		wait for Clk_period;
		Addr <=  "0001011010110";
		Trees_din <= x"b6ff7204";
		wait for Clk_period;
		Addr <=  "0001011010111";
		Trees_din <= x"ff930b89";
		wait for Clk_period;
		Addr <=  "0001011011000";
		Trees_din <= x"16ff1d04";
		wait for Clk_period;
		Addr <=  "0001011011001";
		Trees_din <= x"00380b89";
		wait for Clk_period;
		Addr <=  "0001011011010";
		Trees_din <= x"013f0b89";
		wait for Clk_period;
		Addr <=  "0001011011011";
		Trees_din <= x"cbff6608";
		wait for Clk_period;
		Addr <=  "0001011011100";
		Trees_din <= x"6affcf04";
		wait for Clk_period;
		Addr <=  "0001011011101";
		Trees_din <= x"00090b89";
		wait for Clk_period;
		Addr <=  "0001011011110";
		Trees_din <= x"011c0b89";
		wait for Clk_period;
		Addr <=  "0001011011111";
		Trees_din <= x"32ff8104";
		wait for Clk_period;
		Addr <=  "0001011100000";
		Trees_din <= x"ff8f0b89";
		wait for Clk_period;
		Addr <=  "0001011100001";
		Trees_din <= x"00280b89";
		wait for Clk_period;
		Addr <=  "0001011100010";
		Trees_din <= x"a1ff2838";
		wait for Clk_period;
		Addr <=  "0001011100011";
		Trees_din <= x"7b002d28";
		wait for Clk_period;
		Addr <=  "0001011100100";
		Trees_din <= x"9ffffe18";
		wait for Clk_period;
		Addr <=  "0001011100101";
		Trees_din <= x"a6fe9d08";
		wait for Clk_period;
		Addr <=  "0001011100110";
		Trees_din <= x"64febe04";
		wait for Clk_period;
		Addr <=  "0001011100111";
		Trees_din <= x"00e60cdd";
		wait for Clk_period;
		Addr <=  "0001011101000";
		Trees_din <= x"ff920cdd";
		wait for Clk_period;
		Addr <=  "0001011101001";
		Trees_din <= x"f6fe0c08";
		wait for Clk_period;
		Addr <=  "0001011101010";
		Trees_din <= x"c7feff04";
		wait for Clk_period;
		Addr <=  "0001011101011";
		Trees_din <= x"ffa90cdd";
		wait for Clk_period;
		Addr <=  "0001011101100";
		Trees_din <= x"00a20cdd";
		wait for Clk_period;
		Addr <=  "0001011101101";
		Trees_din <= x"35ffe004";
		wait for Clk_period;
		Addr <=  "0001011101110";
		Trees_din <= x"ff6f0cdd";
		wait for Clk_period;
		Addr <=  "0001011101111";
		Trees_din <= x"000c0cdd";
		wait for Clk_period;
		Addr <=  "0001011110000";
		Trees_din <= x"d4ff8404";
		wait for Clk_period;
		Addr <=  "0001011110001";
		Trees_din <= x"ff880cdd";
		wait for Clk_period;
		Addr <=  "0001011110010";
		Trees_din <= x"68ff1a08";
		wait for Clk_period;
		Addr <=  "0001011110011";
		Trees_din <= x"a4ff9204";
		wait for Clk_period;
		Addr <=  "0001011110100";
		Trees_din <= x"00f00cdd";
		wait for Clk_period;
		Addr <=  "0001011110101";
		Trees_din <= x"00330cdd";
		wait for Clk_period;
		Addr <=  "0001011110110";
		Trees_din <= x"ffe30cdd";
		wait for Clk_period;
		Addr <=  "0001011110111";
		Trees_din <= x"5efff30c";
		wait for Clk_period;
		Addr <=  "0001011111000";
		Trees_din <= x"ba002408";
		wait for Clk_period;
		Addr <=  "0001011111001";
		Trees_din <= x"8effde04";
		wait for Clk_period;
		Addr <=  "0001011111010";
		Trees_din <= x"011a0cdd";
		wait for Clk_period;
		Addr <=  "0001011111011";
		Trees_din <= x"005b0cdd";
		wait for Clk_period;
		Addr <=  "0001011111100";
		Trees_din <= x"fff50cdd";
		wait for Clk_period;
		Addr <=  "0001011111101";
		Trees_din <= x"ff900cdd";
		wait for Clk_period;
		Addr <=  "0001011111110";
		Trees_din <= x"16ff0c38";
		wait for Clk_period;
		Addr <=  "0001011111111";
		Trees_din <= x"d3fe951c";
		wait for Clk_period;
		Addr <=  "0001100000000";
		Trees_din <= x"9dffc510";
		wait for Clk_period;
		Addr <=  "0001100000001";
		Trees_din <= x"41ff7708";
		wait for Clk_period;
		Addr <=  "0001100000010";
		Trees_din <= x"2e001c04";
		wait for Clk_period;
		Addr <=  "0001100000011";
		Trees_din <= x"ff6e0cdd";
		wait for Clk_period;
		Addr <=  "0001100000100";
		Trees_din <= x"002e0cdd";
		wait for Clk_period;
		Addr <=  "0001100000101";
		Trees_din <= x"57ff7d04";
		wait for Clk_period;
		Addr <=  "0001100000110";
		Trees_din <= x"fffb0cdd";
		wait for Clk_period;
		Addr <=  "0001100000111";
		Trees_din <= x"00bc0cdd";
		wait for Clk_period;
		Addr <=  "0001100001000";
		Trees_din <= x"d8003704";
		wait for Clk_period;
		Addr <=  "0001100001001";
		Trees_din <= x"ff9f0cdd";
		wait for Clk_period;
		Addr <=  "0001100001010";
		Trees_din <= x"47000704";
		wait for Clk_period;
		Addr <=  "0001100001011";
		Trees_din <= x"00fb0cdd";
		wait for Clk_period;
		Addr <=  "0001100001100";
		Trees_din <= x"ffd80cdd";
		wait for Clk_period;
		Addr <=  "0001100001101";
		Trees_din <= x"f6fe400c";
		wait for Clk_period;
		Addr <=  "0001100001110";
		Trees_din <= x"19ffb308";
		wait for Clk_period;
		Addr <=  "0001100001111";
		Trees_din <= x"57003b04";
		wait for Clk_period;
		Addr <=  "0001100010000";
		Trees_din <= x"ff8e0cdd";
		wait for Clk_period;
		Addr <=  "0001100010001";
		Trees_din <= x"00620cdd";
		wait for Clk_period;
		Addr <=  "0001100010010";
		Trees_din <= x"00be0cdd";
		wait for Clk_period;
		Addr <=  "0001100010011";
		Trees_din <= x"35ffd908";
		wait for Clk_period;
		Addr <=  "0001100010100";
		Trees_din <= x"8cfe8a04";
		wait for Clk_period;
		Addr <=  "0001100010101";
		Trees_din <= x"00780cdd";
		wait for Clk_period;
		Addr <=  "0001100010110";
		Trees_din <= x"ff700cdd";
		wait for Clk_period;
		Addr <=  "0001100010111";
		Trees_din <= x"c4ff5504";
		wait for Clk_period;
		Addr <=  "0001100011000";
		Trees_din <= x"00790cdd";
		wait for Clk_period;
		Addr <=  "0001100011001";
		Trees_din <= x"ff8c0cdd";
		wait for Clk_period;
		Addr <=  "0001100011010";
		Trees_din <= x"b3ff3b20";
		wait for Clk_period;
		Addr <=  "0001100011011";
		Trees_din <= x"52fee510";
		wait for Clk_period;
		Addr <=  "0001100011100";
		Trees_din <= x"e0feda08";
		wait for Clk_period;
		Addr <=  "0001100011101";
		Trees_din <= x"beffa604";
		wait for Clk_period;
		Addr <=  "0001100011110";
		Trees_din <= x"00ba0cdd";
		wait for Clk_period;
		Addr <=  "0001100011111";
		Trees_din <= x"ff910cdd";
		wait for Clk_period;
		Addr <=  "0001100100000";
		Trees_din <= x"de002604";
		wait for Clk_period;
		Addr <=  "0001100100001";
		Trees_din <= x"ff6c0cdd";
		wait for Clk_period;
		Addr <=  "0001100100010";
		Trees_din <= x"00060cdd";
		wait for Clk_period;
		Addr <=  "0001100100011";
		Trees_din <= x"f8007f08";
		wait for Clk_period;
		Addr <=  "0001100100100";
		Trees_din <= x"ecffa904";
		wait for Clk_period;
		Addr <=  "0001100100101";
		Trees_din <= x"ffec0cdd";
		wait for Clk_period;
		Addr <=  "0001100100110";
		Trees_din <= x"00be0cdd";
		wait for Clk_period;
		Addr <=  "0001100100111";
		Trees_din <= x"6aff0004";
		wait for Clk_period;
		Addr <=  "0001100101000";
		Trees_din <= x"00bf0cdd";
		wait for Clk_period;
		Addr <=  "0001100101001";
		Trees_din <= x"ffbf0cdd";
		wait for Clk_period;
		Addr <=  "0001100101010";
		Trees_din <= x"beff520c";
		wait for Clk_period;
		Addr <=  "0001100101011";
		Trees_din <= x"a2ffcd08";
		wait for Clk_period;
		Addr <=  "0001100101100";
		Trees_din <= x"1aff0904";
		wait for Clk_period;
		Addr <=  "0001100101101";
		Trees_din <= x"00290cdd";
		wait for Clk_period;
		Addr <=  "0001100101110";
		Trees_din <= x"00e00cdd";
		wait for Clk_period;
		Addr <=  "0001100101111";
		Trees_din <= x"ffa70cdd";
		wait for Clk_period;
		Addr <=  "0001100110000";
		Trees_din <= x"f1fffc08";
		wait for Clk_period;
		Addr <=  "0001100110001";
		Trees_din <= x"14007f04";
		wait for Clk_period;
		Addr <=  "0001100110010";
		Trees_din <= x"ff660cdd";
		wait for Clk_period;
		Addr <=  "0001100110011";
		Trees_din <= x"00480cdd";
		wait for Clk_period;
		Addr <=  "0001100110100";
		Trees_din <= x"d9ffd504";
		wait for Clk_period;
		Addr <=  "0001100110101";
		Trees_din <= x"ffa40cdd";
		wait for Clk_period;
		Addr <=  "0001100110110";
		Trees_din <= x"01000cdd";
		wait for Clk_period;
		Addr <=  "0001100110111";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0001100111000";
		Trees_din <= x"2200ac58";
		wait for Clk_period;
		Addr <=  "0001100111001";
		Trees_din <= x"47002534";
		wait for Clk_period;
		Addr <=  "0001100111010";
		Trees_din <= x"41feb914";
		wait for Clk_period;
		Addr <=  "0001100111011";
		Trees_din <= x"a5ffd90c";
		wait for Clk_period;
		Addr <=  "0001100111100";
		Trees_din <= x"57007808";
		wait for Clk_period;
		Addr <=  "0001100111101";
		Trees_din <= x"f6fe0004";
		wait for Clk_period;
		Addr <=  "0001100111110";
		Trees_din <= x"003f0dc5";
		wait for Clk_period;
		Addr <=  "0001100111111";
		Trees_din <= x"ff670dc5";
		wait for Clk_period;
		Addr <=  "0001101000000";
		Trees_din <= x"00690dc5";
		wait for Clk_period;
		Addr <=  "0001101000001";
		Trees_din <= x"41fe4304";
		wait for Clk_period;
		Addr <=  "0001101000010";
		Trees_din <= x"009b0dc5";
		wait for Clk_period;
		Addr <=  "0001101000011";
		Trees_din <= x"001a0dc5";
		wait for Clk_period;
		Addr <=  "0001101000100";
		Trees_din <= x"18000410";
		wait for Clk_period;
		Addr <=  "0001101000101";
		Trees_din <= x"6cff2708";
		wait for Clk_period;
		Addr <=  "0001101000110";
		Trees_din <= x"7affd304";
		wait for Clk_period;
		Addr <=  "0001101000111";
		Trees_din <= x"00b20dc5";
		wait for Clk_period;
		Addr <=  "0001101001000";
		Trees_din <= x"fff60dc5";
		wait for Clk_period;
		Addr <=  "0001101001001";
		Trees_din <= x"68fedd04";
		wait for Clk_period;
		Addr <=  "0001101001010";
		Trees_din <= x"004d0dc5";
		wait for Clk_period;
		Addr <=  "0001101001011";
		Trees_din <= x"ffc70dc5";
		wait for Clk_period;
		Addr <=  "0001101001100";
		Trees_din <= x"02ff2208";
		wait for Clk_period;
		Addr <=  "0001101001101";
		Trees_din <= x"80001704";
		wait for Clk_period;
		Addr <=  "0001101001110";
		Trees_din <= x"ff690dc5";
		wait for Clk_period;
		Addr <=  "0001101001111";
		Trees_din <= x"00350dc5";
		wait for Clk_period;
		Addr <=  "0001101010000";
		Trees_din <= x"3dffb904";
		wait for Clk_period;
		Addr <=  "0001101010001";
		Trees_din <= x"00a00dc5";
		wait for Clk_period;
		Addr <=  "0001101010010";
		Trees_din <= x"ff840dc5";
		wait for Clk_period;
		Addr <=  "0001101010011";
		Trees_din <= x"35ffd910";
		wait for Clk_period;
		Addr <=  "0001101010100";
		Trees_din <= x"a400200c";
		wait for Clk_period;
		Addr <=  "0001101010101";
		Trees_din <= x"d3fe0704";
		wait for Clk_period;
		Addr <=  "0001101010110";
		Trees_din <= x"00710dc5";
		wait for Clk_period;
		Addr <=  "0001101010111";
		Trees_din <= x"16ff8304";
		wait for Clk_period;
		Addr <=  "0001101011000";
		Trees_din <= x"ff700dc5";
		wait for Clk_period;
		Addr <=  "0001101011001";
		Trees_din <= x"ffea0dc5";
		wait for Clk_period;
		Addr <=  "0001101011010";
		Trees_din <= x"00af0dc5";
		wait for Clk_period;
		Addr <=  "0001101011011";
		Trees_din <= x"8fff0604";
		wait for Clk_period;
		Addr <=  "0001101011100";
		Trees_din <= x"ff8c0dc5";
		wait for Clk_period;
		Addr <=  "0001101011101";
		Trees_din <= x"f4fe7408";
		wait for Clk_period;
		Addr <=  "0001101011110";
		Trees_din <= x"0500b004";
		wait for Clk_period;
		Addr <=  "0001101011111";
		Trees_din <= x"ff9d0dc5";
		wait for Clk_period;
		Addr <=  "0001101100000";
		Trees_din <= x"00070dc5";
		wait for Clk_period;
		Addr <=  "0001101100001";
		Trees_din <= x"ebfed304";
		wait for Clk_period;
		Addr <=  "0001101100010";
		Trees_din <= x"fffb0dc5";
		wait for Clk_period;
		Addr <=  "0001101100011";
		Trees_din <= x"00c10dc5";
		wait for Clk_period;
		Addr <=  "0001101100100";
		Trees_din <= x"beff7410";
		wait for Clk_period;
		Addr <=  "0001101100101";
		Trees_din <= x"34ffbe08";
		wait for Clk_period;
		Addr <=  "0001101100110";
		Trees_din <= x"e2fefa04";
		wait for Clk_period;
		Addr <=  "0001101100111";
		Trees_din <= x"00d20dc5";
		wait for Clk_period;
		Addr <=  "0001101101000";
		Trees_din <= x"fffb0dc5";
		wait for Clk_period;
		Addr <=  "0001101101001";
		Trees_din <= x"57ffc104";
		wait for Clk_period;
		Addr <=  "0001101101010";
		Trees_din <= x"ff730dc5";
		wait for Clk_period;
		Addr <=  "0001101101011";
		Trees_din <= x"00470dc5";
		wait for Clk_period;
		Addr <=  "0001101101100";
		Trees_din <= x"a9fe7a08";
		wait for Clk_period;
		Addr <=  "0001101101101";
		Trees_din <= x"01fecb04";
		wait for Clk_period;
		Addr <=  "0001101101110";
		Trees_din <= x"ffb00dc5";
		wait for Clk_period;
		Addr <=  "0001101101111";
		Trees_din <= x"00b70dc5";
		wait for Clk_period;
		Addr <=  "0001101110000";
		Trees_din <= x"ff650dc5";
		wait for Clk_period;
		Addr <=  "0001101110001";
		Trees_din <= x"2200ac40";
		wait for Clk_period;
		Addr <=  "0001101110010";
		Trees_din <= x"23000728";
		wait for Clk_period;
		Addr <=  "0001101110011";
		Trees_din <= x"2a00bb20";
		wait for Clk_period;
		Addr <=  "0001101110100";
		Trees_din <= x"a2ff9910";
		wait for Clk_period;
		Addr <=  "0001101110101";
		Trees_din <= x"36fedd08";
		wait for Clk_period;
		Addr <=  "0001101110110";
		Trees_din <= x"01fe9e04";
		wait for Clk_period;
		Addr <=  "0001101110111";
		Trees_din <= x"ffac0e81";
		wait for Clk_period;
		Addr <=  "0001101111000";
		Trees_din <= x"00b90e81";
		wait for Clk_period;
		Addr <=  "0001101111001";
		Trees_din <= x"cafeea04";
		wait for Clk_period;
		Addr <=  "0001101111010";
		Trees_din <= x"ff7b0e81";
		wait for Clk_period;
		Addr <=  "0001101111011";
		Trees_din <= x"002c0e81";
		wait for Clk_period;
		Addr <=  "0001101111100";
		Trees_din <= x"faff8e08";
		wait for Clk_period;
		Addr <=  "0001101111101";
		Trees_din <= x"18001904";
		wait for Clk_period;
		Addr <=  "0001101111110";
		Trees_din <= x"00660e81";
		wait for Clk_period;
		Addr <=  "0001101111111";
		Trees_din <= x"ffb50e81";
		wait for Clk_period;
		Addr <=  "0001110000000";
		Trees_din <= x"f1001904";
		wait for Clk_period;
		Addr <=  "0001110000001";
		Trees_din <= x"ffb50e81";
		wait for Clk_period;
		Addr <=  "0001110000010";
		Trees_din <= x"005a0e81";
		wait for Clk_period;
		Addr <=  "0001110000011";
		Trees_din <= x"7eff7404";
		wait for Clk_period;
		Addr <=  "0001110000100";
		Trees_din <= x"ff6a0e81";
		wait for Clk_period;
		Addr <=  "0001110000101";
		Trees_din <= x"003e0e81";
		wait for Clk_period;
		Addr <=  "0001110000110";
		Trees_din <= x"49fef308";
		wait for Clk_period;
		Addr <=  "0001110000111";
		Trees_din <= x"76001904";
		wait for Clk_period;
		Addr <=  "0001110001000";
		Trees_din <= x"ffd90e81";
		wait for Clk_period;
		Addr <=  "0001110001001";
		Trees_din <= x"00b60e81";
		wait for Clk_period;
		Addr <=  "0001110001010";
		Trees_din <= x"f6fe0c04";
		wait for Clk_period;
		Addr <=  "0001110001011";
		Trees_din <= x"00280e81";
		wait for Clk_period;
		Addr <=  "0001110001100";
		Trees_din <= x"9f003108";
		wait for Clk_period;
		Addr <=  "0001110001101";
		Trees_din <= x"ce006404";
		wait for Clk_period;
		Addr <=  "0001110001110";
		Trees_din <= x"ff660e81";
		wait for Clk_period;
		Addr <=  "0001110001111";
		Trees_din <= x"fff30e81";
		wait for Clk_period;
		Addr <=  "0001110010000";
		Trees_din <= x"00120e81";
		wait for Clk_period;
		Addr <=  "0001110010001";
		Trees_din <= x"beff7414";
		wait for Clk_period;
		Addr <=  "0001110010010";
		Trees_din <= x"c7ff4108";
		wait for Clk_period;
		Addr <=  "0001110010011";
		Trees_din <= x"abfff804";
		wait for Clk_period;
		Addr <=  "0001110010100";
		Trees_din <= x"002c0e81";
		wait for Clk_period;
		Addr <=  "0001110010101";
		Trees_din <= x"ff770e81";
		wait for Clk_period;
		Addr <=  "0001110010110";
		Trees_din <= x"83ff1f08";
		wait for Clk_period;
		Addr <=  "0001110010111";
		Trees_din <= x"b1ff3504";
		wait for Clk_period;
		Addr <=  "0001110011000";
		Trees_din <= x"00260e81";
		wait for Clk_period;
		Addr <=  "0001110011001";
		Trees_din <= x"00c60e81";
		wait for Clk_period;
		Addr <=  "0001110011010";
		Trees_din <= x"ffaa0e81";
		wait for Clk_period;
		Addr <=  "0001110011011";
		Trees_din <= x"a9fe7a08";
		wait for Clk_period;
		Addr <=  "0001110011100";
		Trees_din <= x"05008704";
		wait for Clk_period;
		Addr <=  "0001110011101";
		Trees_din <= x"ffb10e81";
		wait for Clk_period;
		Addr <=  "0001110011110";
		Trees_din <= x"00ac0e81";
		wait for Clk_period;
		Addr <=  "0001110011111";
		Trees_din <= x"ff660e81";
		wait for Clk_period;
		Addr <=  "0001110100000";
		Trees_din <= x"f202686c";
		wait for Clk_period;
		Addr <=  "0001110100001";
		Trees_din <= x"6cff643c";
		wait for Clk_period;
		Addr <=  "0001110100010";
		Trees_din <= x"d2feb620";
		wait for Clk_period;
		Addr <=  "0001110100011";
		Trees_din <= x"9bfec410";
		wait for Clk_period;
		Addr <=  "0001110100100";
		Trees_din <= x"87ff5308";
		wait for Clk_period;
		Addr <=  "0001110100101";
		Trees_din <= x"baff4504";
		wait for Clk_period;
		Addr <=  "0001110100110";
		Trees_din <= x"004c0fbd";
		wait for Clk_period;
		Addr <=  "0001110100111";
		Trees_din <= x"ff860fbd";
		wait for Clk_period;
		Addr <=  "0001110101000";
		Trees_din <= x"81ff7904";
		wait for Clk_period;
		Addr <=  "0001110101001";
		Trees_din <= x"00c10fbd";
		wait for Clk_period;
		Addr <=  "0001110101010";
		Trees_din <= x"ffac0fbd";
		wait for Clk_period;
		Addr <=  "0001110101011";
		Trees_din <= x"61fef608";
		wait for Clk_period;
		Addr <=  "0001110101100";
		Trees_din <= x"01feee04";
		wait for Clk_period;
		Addr <=  "0001110101101";
		Trees_din <= x"ff900fbd";
		wait for Clk_period;
		Addr <=  "0001110101110";
		Trees_din <= x"00790fbd";
		wait for Clk_period;
		Addr <=  "0001110101111";
		Trees_din <= x"afff1904";
		wait for Clk_period;
		Addr <=  "0001110110000";
		Trees_din <= x"002b0fbd";
		wait for Clk_period;
		Addr <=  "0001110110001";
		Trees_din <= x"ff690fbd";
		wait for Clk_period;
		Addr <=  "0001110110010";
		Trees_din <= x"f0ff930c";
		wait for Clk_period;
		Addr <=  "0001110110011";
		Trees_din <= x"70ffa208";
		wait for Clk_period;
		Addr <=  "0001110110100";
		Trees_din <= x"4afed504";
		wait for Clk_period;
		Addr <=  "0001110110101";
		Trees_din <= x"ffd70fbd";
		wait for Clk_period;
		Addr <=  "0001110110110";
		Trees_din <= x"00820fbd";
		wait for Clk_period;
		Addr <=  "0001110110111";
		Trees_din <= x"ff840fbd";
		wait for Clk_period;
		Addr <=  "0001110111000";
		Trees_din <= x"3afec208";
		wait for Clk_period;
		Addr <=  "0001110111001";
		Trees_din <= x"f5000504";
		wait for Clk_period;
		Addr <=  "0001110111010";
		Trees_din <= x"00cb0fbd";
		wait for Clk_period;
		Addr <=  "0001110111011";
		Trees_din <= x"fff20fbd";
		wait for Clk_period;
		Addr <=  "0001110111100";
		Trees_din <= x"0efe2104";
		wait for Clk_period;
		Addr <=  "0001110111101";
		Trees_din <= x"00950fbd";
		wait for Clk_period;
		Addr <=  "0001110111110";
		Trees_din <= x"ff880fbd";
		wait for Clk_period;
		Addr <=  "0001110111111";
		Trees_din <= x"6ffeeb10";
		wait for Clk_period;
		Addr <=  "0001111000000";
		Trees_din <= x"dcff9e04";
		wait for Clk_period;
		Addr <=  "0001111000001";
		Trees_din <= x"ff8b0fbd";
		wait for Clk_period;
		Addr <=  "0001111000010";
		Trees_din <= x"4fffb108";
		wait for Clk_period;
		Addr <=  "0001111000011";
		Trees_din <= x"4eff6c04";
		wait for Clk_period;
		Addr <=  "0001111000100";
		Trees_din <= x"00070fbd";
		wait for Clk_period;
		Addr <=  "0001111000101";
		Trees_din <= x"00ec0fbd";
		wait for Clk_period;
		Addr <=  "0001111000110";
		Trees_din <= x"ffd60fbd";
		wait for Clk_period;
		Addr <=  "0001111000111";
		Trees_din <= x"c5ff4b10";
		wait for Clk_period;
		Addr <=  "0001111001000";
		Trees_din <= x"3afe9608";
		wait for Clk_period;
		Addr <=  "0001111001001";
		Trees_din <= x"95ff7104";
		wait for Clk_period;
		Addr <=  "0001111001010";
		Trees_din <= x"ffcf0fbd";
		wait for Clk_period;
		Addr <=  "0001111001011";
		Trees_din <= x"00840fbd";
		wait for Clk_period;
		Addr <=  "0001111001100";
		Trees_din <= x"35002304";
		wait for Clk_period;
		Addr <=  "0001111001101";
		Trees_din <= x"ff660fbd";
		wait for Clk_period;
		Addr <=  "0001111001110";
		Trees_din <= x"00230fbd";
		wait for Clk_period;
		Addr <=  "0001111001111";
		Trees_din <= x"eefffd08";
		wait for Clk_period;
		Addr <=  "0001111010000";
		Trees_din <= x"e5fec504";
		wait for Clk_period;
		Addr <=  "0001111010001";
		Trees_din <= x"00530fbd";
		wait for Clk_period;
		Addr <=  "0001111010010";
		Trees_din <= x"ffa50fbd";
		wait for Clk_period;
		Addr <=  "0001111010011";
		Trees_din <= x"cfff5504";
		wait for Clk_period;
		Addr <=  "0001111010100";
		Trees_din <= x"005f0fbd";
		wait for Clk_period;
		Addr <=  "0001111010101";
		Trees_din <= x"ff770fbd";
		wait for Clk_period;
		Addr <=  "0001111010110";
		Trees_din <= x"a1ff6010";
		wait for Clk_period;
		Addr <=  "0001111010111";
		Trees_din <= x"9a00930c";
		wait for Clk_period;
		Addr <=  "0001111011000";
		Trees_din <= x"8400d708";
		wait for Clk_period;
		Addr <=  "0001111011001";
		Trees_din <= x"f4ffed04";
		wait for Clk_period;
		Addr <=  "0001111011010";
		Trees_din <= x"ff670fbd";
		wait for Clk_period;
		Addr <=  "0001111011011";
		Trees_din <= x"ffeb0fbd";
		wait for Clk_period;
		Addr <=  "0001111011100";
		Trees_din <= x"fff50fbd";
		wait for Clk_period;
		Addr <=  "0001111011101";
		Trees_din <= x"003c0fbd";
		wait for Clk_period;
		Addr <=  "0001111011110";
		Trees_din <= x"3aff2318";
		wait for Clk_period;
		Addr <=  "0001111011111";
		Trees_din <= x"16ff1d0c";
		wait for Clk_period;
		Addr <=  "0001111100000";
		Trees_din <= x"f700d604";
		wait for Clk_period;
		Addr <=  "0001111100001";
		Trees_din <= x"ff7c0fbd";
		wait for Clk_period;
		Addr <=  "0001111100010";
		Trees_din <= x"a7ffc004";
		wait for Clk_period;
		Addr <=  "0001111100011";
		Trees_din <= x"fff90fbd";
		wait for Clk_period;
		Addr <=  "0001111100100";
		Trees_din <= x"00720fbd";
		wait for Clk_period;
		Addr <=  "0001111100101";
		Trees_din <= x"40001404";
		wait for Clk_period;
		Addr <=  "0001111100110";
		Trees_din <= x"ffa60fbd";
		wait for Clk_period;
		Addr <=  "0001111100111";
		Trees_din <= x"2dfeb904";
		wait for Clk_period;
		Addr <=  "0001111101000";
		Trees_din <= x"00ef0fbd";
		wait for Clk_period;
		Addr <=  "0001111101001";
		Trees_din <= x"001e0fbd";
		wait for Clk_period;
		Addr <=  "0001111101010";
		Trees_din <= x"79ffe408";
		wait for Clk_period;
		Addr <=  "0001111101011";
		Trees_din <= x"65feb904";
		wait for Clk_period;
		Addr <=  "0001111101100";
		Trees_din <= x"ffee0fbd";
		wait for Clk_period;
		Addr <=  "0001111101101";
		Trees_din <= x"ff720fbd";
		wait for Clk_period;
		Addr <=  "0001111101110";
		Trees_din <= x"00630fbd";
		wait for Clk_period;
		Addr <=  "0001111101111";
		Trees_din <= x"16ff1344";
		wait for Clk_period;
		Addr <=  "0001111110000";
		Trees_din <= x"d3fe9520";
		wait for Clk_period;
		Addr <=  "0001111110001";
		Trees_din <= x"96ff5410";
		wait for Clk_period;
		Addr <=  "0001111110010";
		Trees_din <= x"35ffe008";
		wait for Clk_period;
		Addr <=  "0001111110011";
		Trees_din <= x"97ff9504";
		wait for Clk_period;
		Addr <=  "0001111110100";
		Trees_din <= x"ff7610b9";
		wait for Clk_period;
		Addr <=  "0001111110101";
		Trees_din <= x"ffff10b9";
		wait for Clk_period;
		Addr <=  "0001111110110";
		Trees_din <= x"0efdc304";
		wait for Clk_period;
		Addr <=  "0001111110111";
		Trees_din <= x"008010b9";
		wait for Clk_period;
		Addr <=  "0001111111000";
		Trees_din <= x"000610b9";
		wait for Clk_period;
		Addr <=  "0001111111001";
		Trees_din <= x"5bff880c";
		wait for Clk_period;
		Addr <=  "0001111111010";
		Trees_din <= x"3dff8604";
		wait for Clk_period;
		Addr <=  "0001111111011";
		Trees_din <= x"ffa310b9";
		wait for Clk_period;
		Addr <=  "0001111111100";
		Trees_din <= x"d8003804";
		wait for Clk_period;
		Addr <=  "0001111111101";
		Trees_din <= x"ffd610b9";
		wait for Clk_period;
		Addr <=  "0001111111110";
		Trees_din <= x"00bb10b9";
		wait for Clk_period;
		Addr <=  "0001111111111";
		Trees_din <= x"ff8610b9";
		wait for Clk_period;
		Addr <=  "0010000000000";
		Trees_din <= x"aa004c1c";
		wait for Clk_period;
		Addr <=  "0010000000001";
		Trees_din <= x"befeed0c";
		wait for Clk_period;
		Addr <=  "0010000000010";
		Trees_din <= x"b1ff0508";
		wait for Clk_period;
		Addr <=  "0010000000011";
		Trees_din <= x"40003e04";
		wait for Clk_period;
		Addr <=  "0010000000100";
		Trees_din <= x"002410b9";
		wait for Clk_period;
		Addr <=  "0010000000101";
		Trees_din <= x"008b10b9";
		wait for Clk_period;
		Addr <=  "0010000000110";
		Trees_din <= x"ffa410b9";
		wait for Clk_period;
		Addr <=  "0010000000111";
		Trees_din <= x"2e006b08";
		wait for Clk_period;
		Addr <=  "0010000001000";
		Trees_din <= x"57003b04";
		wait for Clk_period;
		Addr <=  "0010000001001";
		Trees_din <= x"ff7c10b9";
		wait for Clk_period;
		Addr <=  "0010000001010";
		Trees_din <= x"004210b9";
		wait for Clk_period;
		Addr <=  "0010000001011";
		Trees_din <= x"38feb604";
		wait for Clk_period;
		Addr <=  "0010000001100";
		Trees_din <= x"00c910b9";
		wait for Clk_period;
		Addr <=  "0010000001101";
		Trees_din <= x"ffcd10b9";
		wait for Clk_period;
		Addr <=  "0010000001110";
		Trees_din <= x"96ffe004";
		wait for Clk_period;
		Addr <=  "0010000001111";
		Trees_din <= x"001710b9";
		wait for Clk_period;
		Addr <=  "0010000010000";
		Trees_din <= x"009610b9";
		wait for Clk_period;
		Addr <=  "0010000010001";
		Trees_din <= x"b9fedb10";
		wait for Clk_period;
		Addr <=  "0010000010010";
		Trees_din <= x"57ffcb0c";
		wait for Clk_period;
		Addr <=  "0010000010011";
		Trees_din <= x"44008c04";
		wait for Clk_period;
		Addr <=  "0010000010100";
		Trees_din <= x"ff6f10b9";
		wait for Clk_period;
		Addr <=  "0010000010101";
		Trees_din <= x"a3fff204";
		wait for Clk_period;
		Addr <=  "0010000010110";
		Trees_din <= x"ffa110b9";
		wait for Clk_period;
		Addr <=  "0010000010111";
		Trees_din <= x"008010b9";
		wait for Clk_period;
		Addr <=  "0010000011000";
		Trees_din <= x"006c10b9";
		wait for Clk_period;
		Addr <=  "0010000011001";
		Trees_din <= x"6fff8a14";
		wait for Clk_period;
		Addr <=  "0010000011010";
		Trees_din <= x"2a00ae0c";
		wait for Clk_period;
		Addr <=  "0010000011011";
		Trees_din <= x"3bffb408";
		wait for Clk_period;
		Addr <=  "0010000011100";
		Trees_din <= x"41fead04";
		wait for Clk_period;
		Addr <=  "0010000011101";
		Trees_din <= x"ffaf10b9";
		wait for Clk_period;
		Addr <=  "0010000011110";
		Trees_din <= x"007a10b9";
		wait for Clk_period;
		Addr <=  "0010000011111";
		Trees_din <= x"ff8810b9";
		wait for Clk_period;
		Addr <=  "0010000100000";
		Trees_din <= x"53ffa804";
		wait for Clk_period;
		Addr <=  "0010000100001";
		Trees_din <= x"ff8010b9";
		wait for Clk_period;
		Addr <=  "0010000100010";
		Trees_din <= x"002210b9";
		wait for Clk_period;
		Addr <=  "0010000100011";
		Trees_din <= x"33ffe610";
		wait for Clk_period;
		Addr <=  "0010000100100";
		Trees_din <= x"acfff808";
		wait for Clk_period;
		Addr <=  "0010000100101";
		Trees_din <= x"83ff1a04";
		wait for Clk_period;
		Addr <=  "0010000100110";
		Trees_din <= x"007d10b9";
		wait for Clk_period;
		Addr <=  "0010000100111";
		Trees_din <= x"ffda10b9";
		wait for Clk_period;
		Addr <=  "0010000101000";
		Trees_din <= x"f6fea504";
		wait for Clk_period;
		Addr <=  "0010000101001";
		Trees_din <= x"000f10b9";
		wait for Clk_period;
		Addr <=  "0010000101010";
		Trees_din <= x"ff7e10b9";
		wait for Clk_period;
		Addr <=  "0010000101011";
		Trees_din <= x"c4ff0304";
		wait for Clk_period;
		Addr <=  "0010000101100";
		Trees_din <= x"00ed10b9";
		wait for Clk_period;
		Addr <=  "0010000101101";
		Trees_din <= x"ffd010b9";
		wait for Clk_period;
		Addr <=  "0010000101110";
		Trees_din <= x"2200b240";
		wait for Clk_period;
		Addr <=  "0010000101111";
		Trees_din <= x"23000728";
		wait for Clk_period;
		Addr <=  "0010000110000";
		Trees_din <= x"2a00bb20";
		wait for Clk_period;
		Addr <=  "0010000110001";
		Trees_din <= x"cbff8710";
		wait for Clk_period;
		Addr <=  "0010000110010";
		Trees_din <= x"81ff4f08";
		wait for Clk_period;
		Addr <=  "0010000110011";
		Trees_din <= x"f5ff9804";
		wait for Clk_period;
		Addr <=  "0010000110100";
		Trees_din <= x"ffc7115d";
		wait for Clk_period;
		Addr <=  "0010000110101";
		Trees_din <= x"00a9115d";
		wait for Clk_period;
		Addr <=  "0010000110110";
		Trees_din <= x"d2fe9c04";
		wait for Clk_period;
		Addr <=  "0010000110111";
		Trees_din <= x"ff93115d";
		wait for Clk_period;
		Addr <=  "0010000111000";
		Trees_din <= x"0041115d";
		wait for Clk_period;
		Addr <=  "0010000111001";
		Trees_din <= x"d2feb908";
		wait for Clk_period;
		Addr <=  "0010000111010";
		Trees_din <= x"f7010f04";
		wait for Clk_period;
		Addr <=  "0010000111011";
		Trees_din <= x"ff95115d";
		wait for Clk_period;
		Addr <=  "0010000111100";
		Trees_din <= x"005f115d";
		wait for Clk_period;
		Addr <=  "0010000111101";
		Trees_din <= x"f6fe6804";
		wait for Clk_period;
		Addr <=  "0010000111110";
		Trees_din <= x"0080115d";
		wait for Clk_period;
		Addr <=  "0010000111111";
		Trees_din <= x"0001115d";
		wait for Clk_period;
		Addr <=  "0010001000000";
		Trees_din <= x"7eff7404";
		wait for Clk_period;
		Addr <=  "0010001000001";
		Trees_din <= x"ff6f115d";
		wait for Clk_period;
		Addr <=  "0010001000010";
		Trees_din <= x"003d115d";
		wait for Clk_period;
		Addr <=  "0010001000011";
		Trees_din <= x"49fef308";
		wait for Clk_period;
		Addr <=  "0010001000100";
		Trees_din <= x"eeffc004";
		wait for Clk_period;
		Addr <=  "0010001000101";
		Trees_din <= x"008d115d";
		wait for Clk_period;
		Addr <=  "0010001000110";
		Trees_din <= x"ffe8115d";
		wait for Clk_period;
		Addr <=  "0010001000111";
		Trees_din <= x"f6fe0c04";
		wait for Clk_period;
		Addr <=  "0010001001000";
		Trees_din <= x"0022115d";
		wait for Clk_period;
		Addr <=  "0010001001001";
		Trees_din <= x"ce006408";
		wait for Clk_period;
		Addr <=  "0010001001010";
		Trees_din <= x"cc008404";
		wait for Clk_period;
		Addr <=  "0010001001011";
		Trees_din <= x"ff6c115d";
		wait for Clk_period;
		Addr <=  "0010001001100";
		Trees_din <= x"ffe7115d";
		wait for Clk_period;
		Addr <=  "0010001001101";
		Trees_din <= x"fff8115d";
		wait for Clk_period;
		Addr <=  "0010001001110";
		Trees_din <= x"91003210";
		wait for Clk_period;
		Addr <=  "0010001001111";
		Trees_din <= x"38fe6904";
		wait for Clk_period;
		Addr <=  "0010001010000";
		Trees_din <= x"0030115d";
		wait for Clk_period;
		Addr <=  "0010001010001";
		Trees_din <= x"fcffc708";
		wait for Clk_period;
		Addr <=  "0010001010010";
		Trees_din <= x"6bfe0b04";
		wait for Clk_period;
		Addr <=  "0010001010011";
		Trees_din <= x"ffe7115d";
		wait for Clk_period;
		Addr <=  "0010001010100";
		Trees_din <= x"ff68115d";
		wait for Clk_period;
		Addr <=  "0010001010101";
		Trees_din <= x"0027115d";
		wait for Clk_period;
		Addr <=  "0010001010110";
		Trees_din <= x"004d115d";
		wait for Clk_period;
		Addr <=  "0010001010111";
		Trees_din <= x"8dfe4b14";
		wait for Clk_period;
		Addr <=  "0010001011000";
		Trees_din <= x"7b002d0c";
		wait for Clk_period;
		Addr <=  "0010001011001";
		Trees_din <= x"ea001108";
		wait for Clk_period;
		Addr <=  "0010001011010";
		Trees_din <= x"69fe5404";
		wait for Clk_period;
		Addr <=  "0010001011011";
		Trees_din <= x"ffff1239";
		wait for Clk_period;
		Addr <=  "0010001011100";
		Trees_din <= x"ff691239";
		wait for Clk_period;
		Addr <=  "0010001011101";
		Trees_din <= x"00291239";
		wait for Clk_period;
		Addr <=  "0010001011110";
		Trees_din <= x"16ff1b04";
		wait for Clk_period;
		Addr <=  "0010001011111";
		Trees_din <= x"ffac1239";
		wait for Clk_period;
		Addr <=  "0010001100000";
		Trees_din <= x"00861239";
		wait for Clk_period;
		Addr <=  "0010001100001";
		Trees_din <= x"16feb220";
		wait for Clk_period;
		Addr <=  "0010001100010";
		Trees_din <= x"a0ff540c";
		wait for Clk_period;
		Addr <=  "0010001100011";
		Trees_din <= x"35fff908";
		wait for Clk_period;
		Addr <=  "0010001100100";
		Trees_din <= x"3cfe8504";
		wait for Clk_period;
		Addr <=  "0010001100101";
		Trees_din <= x"fff01239";
		wait for Clk_period;
		Addr <=  "0010001100110";
		Trees_din <= x"ff6c1239";
		wait for Clk_period;
		Addr <=  "0010001100111";
		Trees_din <= x"00271239";
		wait for Clk_period;
		Addr <=  "0010001101000";
		Trees_din <= x"3afeda08";
		wait for Clk_period;
		Addr <=  "0010001101001";
		Trees_din <= x"91ff5904";
		wait for Clk_period;
		Addr <=  "0010001101010";
		Trees_din <= x"008f1239";
		wait for Clk_period;
		Addr <=  "0010001101011";
		Trees_din <= x"fff71239";
		wait for Clk_period;
		Addr <=  "0010001101100";
		Trees_din <= x"95ffd808";
		wait for Clk_period;
		Addr <=  "0010001101101";
		Trees_din <= x"64febc04";
		wait for Clk_period;
		Addr <=  "0010001101110";
		Trees_din <= x"ffdf1239";
		wait for Clk_period;
		Addr <=  "0010001101111";
		Trees_din <= x"ff7e1239";
		wait for Clk_period;
		Addr <=  "0010001110000";
		Trees_din <= x"005a1239";
		wait for Clk_period;
		Addr <=  "0010001110001";
		Trees_din <= x"18000420";
		wait for Clk_period;
		Addr <=  "0010001110010";
		Trees_din <= x"47004410";
		wait for Clk_period;
		Addr <=  "0010001110011";
		Trees_din <= x"a2ff9908";
		wait for Clk_period;
		Addr <=  "0010001110100";
		Trees_din <= x"afff6704";
		wait for Clk_period;
		Addr <=  "0010001110101";
		Trees_din <= x"00361239";
		wait for Clk_period;
		Addr <=  "0010001110110";
		Trees_din <= x"ff901239";
		wait for Clk_period;
		Addr <=  "0010001110111";
		Trees_din <= x"faff8d04";
		wait for Clk_period;
		Addr <=  "0010001111000";
		Trees_din <= x"00601239";
		wait for Clk_period;
		Addr <=  "0010001111001";
		Trees_din <= x"fffa1239";
		wait for Clk_period;
		Addr <=  "0010001111010";
		Trees_din <= x"f1000308";
		wait for Clk_period;
		Addr <=  "0010001111011";
		Trees_din <= x"fb006004";
		wait for Clk_period;
		Addr <=  "0010001111100";
		Trees_din <= x"ff711239";
		wait for Clk_period;
		Addr <=  "0010001111101";
		Trees_din <= x"00241239";
		wait for Clk_period;
		Addr <=  "0010001111110";
		Trees_din <= x"78ff9a04";
		wait for Clk_period;
		Addr <=  "0010001111111";
		Trees_din <= x"ffc91239";
		wait for Clk_period;
		Addr <=  "0010010000000";
		Trees_din <= x"00831239";
		wait for Clk_period;
		Addr <=  "0010010000001";
		Trees_din <= x"02ff1d0c";
		wait for Clk_period;
		Addr <=  "0010010000010";
		Trees_din <= x"0ffe9f04";
		wait for Clk_period;
		Addr <=  "0010010000011";
		Trees_din <= x"004f1239";
		wait for Clk_period;
		Addr <=  "0010010000100";
		Trees_din <= x"6ffeeb04";
		wait for Clk_period;
		Addr <=  "0010010000101";
		Trees_din <= x"00041239";
		wait for Clk_period;
		Addr <=  "0010010000110";
		Trees_din <= x"ff6c1239";
		wait for Clk_period;
		Addr <=  "0010010000111";
		Trees_din <= x"4bff0108";
		wait for Clk_period;
		Addr <=  "0010010001000";
		Trees_din <= x"54003104";
		wait for Clk_period;
		Addr <=  "0010010001001";
		Trees_din <= x"ffb11239";
		wait for Clk_period;
		Addr <=  "0010010001010";
		Trees_din <= x"009c1239";
		wait for Clk_period;
		Addr <=  "0010010001011";
		Trees_din <= x"50ff6804";
		wait for Clk_period;
		Addr <=  "0010010001100";
		Trees_din <= x"ff911239";
		wait for Clk_period;
		Addr <=  "0010010001101";
		Trees_din <= x"fffc1239";
		wait for Clk_period;
		Addr <=  "0010010001110";
		Trees_din <= x"16ff0c38";
		wait for Clk_period;
		Addr <=  "0010010001111";
		Trees_din <= x"d3fe9518";
		wait for Clk_period;
		Addr <=  "0010010010000";
		Trees_din <= x"6cffbc14";
		wait for Clk_period;
		Addr <=  "0010010010001";
		Trees_din <= x"d8003808";
		wait for Clk_period;
		Addr <=  "0010010010010";
		Trees_din <= x"32fe6304";
		wait for Clk_period;
		Addr <=  "0010010010011";
		Trees_din <= x"0036131d";
		wait for Clk_period;
		Addr <=  "0010010010100";
		Trees_din <= x"ff88131d";
		wait for Clk_period;
		Addr <=  "0010010010101";
		Trees_din <= x"3dff8604";
		wait for Clk_period;
		Addr <=  "0010010010110";
		Trees_din <= x"ffa8131d";
		wait for Clk_period;
		Addr <=  "0010010010111";
		Trees_din <= x"96ff3904";
		wait for Clk_period;
		Addr <=  "0010010011000";
		Trees_din <= x"ffbc131d";
		wait for Clk_period;
		Addr <=  "0010010011001";
		Trees_din <= x"0090131d";
		wait for Clk_period;
		Addr <=  "0010010011010";
		Trees_din <= x"ff87131d";
		wait for Clk_period;
		Addr <=  "0010010011011";
		Trees_din <= x"57003b18";
		wait for Clk_period;
		Addr <=  "0010010011100";
		Trees_din <= x"96001d10";
		wait for Clk_period;
		Addr <=  "0010010011101";
		Trees_din <= x"35ffd908";
		wait for Clk_period;
		Addr <=  "0010010011110";
		Trees_din <= x"f6fe4004";
		wait for Clk_period;
		Addr <=  "0010010011111";
		Trees_din <= x"fffb131d";
		wait for Clk_period;
		Addr <=  "0010010100000";
		Trees_din <= x"ff72131d";
		wait for Clk_period;
		Addr <=  "0010010100001";
		Trees_din <= x"c4ff5504";
		wait for Clk_period;
		Addr <=  "0010010100010";
		Trees_din <= x"006d131d";
		wait for Clk_period;
		Addr <=  "0010010100011";
		Trees_din <= x"ff97131d";
		wait for Clk_period;
		Addr <=  "0010010100100";
		Trees_din <= x"8cff0204";
		wait for Clk_period;
		Addr <=  "0010010100101";
		Trees_din <= x"009d131d";
		wait for Clk_period;
		Addr <=  "0010010100110";
		Trees_din <= x"ffb0131d";
		wait for Clk_period;
		Addr <=  "0010010100111";
		Trees_din <= x"91ff5804";
		wait for Clk_period;
		Addr <=  "0010010101000";
		Trees_din <= x"0075131d";
		wait for Clk_period;
		Addr <=  "0010010101001";
		Trees_din <= x"0016131d";
		wait for Clk_period;
		Addr <=  "0010010101010";
		Trees_din <= x"b9fedb10";
		wait for Clk_period;
		Addr <=  "0010010101011";
		Trees_din <= x"15fefb04";
		wait for Clk_period;
		Addr <=  "0010010101100";
		Trees_din <= x"0051131d";
		wait for Clk_period;
		Addr <=  "0010010101101";
		Trees_din <= x"55ff8208";
		wait for Clk_period;
		Addr <=  "0010010101110";
		Trees_din <= x"9bfee404";
		wait for Clk_period;
		Addr <=  "0010010101111";
		Trees_din <= x"005a131d";
		wait for Clk_period;
		Addr <=  "0010010110000";
		Trees_din <= x"ffce131d";
		wait for Clk_period;
		Addr <=  "0010010110001";
		Trees_din <= x"ff6f131d";
		wait for Clk_period;
		Addr <=  "0010010110010";
		Trees_din <= x"83ff3a10";
		wait for Clk_period;
		Addr <=  "0010010110011";
		Trees_din <= x"61ffda0c";
		wait for Clk_period;
		Addr <=  "0010010110100";
		Trees_din <= x"c4ffd108";
		wait for Clk_period;
		Addr <=  "0010010110101";
		Trees_din <= x"34001f04";
		wait for Clk_period;
		Addr <=  "0010010110110";
		Trees_din <= x"0078131d";
		wait for Clk_period;
		Addr <=  "0010010110111";
		Trees_din <= x"fffb131d";
		wait for Clk_period;
		Addr <=  "0010010111000";
		Trees_din <= x"ffa3131d";
		wait for Clk_period;
		Addr <=  "0010010111001";
		Trees_din <= x"ff80131d";
		wait for Clk_period;
		Addr <=  "0010010111010";
		Trees_din <= x"85ffce0c";
		wait for Clk_period;
		Addr <=  "0010010111011";
		Trees_din <= x"4400ad08";
		wait for Clk_period;
		Addr <=  "0010010111100";
		Trees_din <= x"3effde04";
		wait for Clk_period;
		Addr <=  "0010010111101";
		Trees_din <= x"ff91131d";
		wait for Clk_period;
		Addr <=  "0010010111110";
		Trees_din <= x"006c131d";
		wait for Clk_period;
		Addr <=  "0010010111111";
		Trees_din <= x"00a5131d";
		wait for Clk_period;
		Addr <=  "0010011000000";
		Trees_din <= x"46ff3d08";
		wait for Clk_period;
		Addr <=  "0010011000001";
		Trees_din <= x"adffb804";
		wait for Clk_period;
		Addr <=  "0010011000010";
		Trees_din <= x"ff88131d";
		wait for Clk_period;
		Addr <=  "0010011000011";
		Trees_din <= x"0043131d";
		wait for Clk_period;
		Addr <=  "0010011000100";
		Trees_din <= x"2bffd704";
		wait for Clk_period;
		Addr <=  "0010011000101";
		Trees_din <= x"008f131d";
		wait for Clk_period;
		Addr <=  "0010011000110";
		Trees_din <= x"ffb5131d";
		wait for Clk_period;
		Addr <=  "0010011000111";
		Trees_din <= x"2200ac48";
		wait for Clk_period;
		Addr <=  "0010011001000";
		Trees_din <= x"2a00a13c";
		wait for Clk_period;
		Addr <=  "0010011001001";
		Trees_din <= x"cbffce1c";
		wait for Clk_period;
		Addr <=  "0010011001010";
		Trees_din <= x"41feb90c";
		wait for Clk_period;
		Addr <=  "0010011001011";
		Trees_din <= x"57007808";
		wait for Clk_period;
		Addr <=  "0010011001100";
		Trees_din <= x"06fee504";
		wait for Clk_period;
		Addr <=  "0010011001101";
		Trees_din <= x"002713d9";
		wait for Clk_period;
		Addr <=  "0010011001110";
		Trees_din <= x"ff8313d9";
		wait for Clk_period;
		Addr <=  "0010011001111";
		Trees_din <= x"006e13d9";
		wait for Clk_period;
		Addr <=  "0010011010000";
		Trees_din <= x"b3ff4b08";
		wait for Clk_period;
		Addr <=  "0010011010001";
		Trees_din <= x"c1fedf04";
		wait for Clk_period;
		Addr <=  "0010011010010";
		Trees_din <= x"006213d9";
		wait for Clk_period;
		Addr <=  "0010011010011";
		Trees_din <= x"000313d9";
		wait for Clk_period;
		Addr <=  "0010011010100";
		Trees_din <= x"18ff6204";
		wait for Clk_period;
		Addr <=  "0010011010101";
		Trees_din <= x"004013d9";
		wait for Clk_period;
		Addr <=  "0010011010110";
		Trees_din <= x"ff9e13d9";
		wait for Clk_period;
		Addr <=  "0010011010111";
		Trees_din <= x"c4fee010";
		wait for Clk_period;
		Addr <=  "0010011011000";
		Trees_din <= x"b4ff1508";
		wait for Clk_period;
		Addr <=  "0010011011001";
		Trees_din <= x"89005204";
		wait for Clk_period;
		Addr <=  "0010011011010";
		Trees_din <= x"ff9313d9";
		wait for Clk_period;
		Addr <=  "0010011011011";
		Trees_din <= x"003813d9";
		wait for Clk_period;
		Addr <=  "0010011011100";
		Trees_din <= x"d2feb504";
		wait for Clk_period;
		Addr <=  "0010011011101";
		Trees_din <= x"ffab13d9";
		wait for Clk_period;
		Addr <=  "0010011011110";
		Trees_din <= x"009513d9";
		wait for Clk_period;
		Addr <=  "0010011011111";
		Trees_din <= x"d600e308";
		wait for Clk_period;
		Addr <=  "0010011100000";
		Trees_din <= x"3dff4004";
		wait for Clk_period;
		Addr <=  "0010011100001";
		Trees_din <= x"004613d9";
		wait for Clk_period;
		Addr <=  "0010011100010";
		Trees_din <= x"ff8a13d9";
		wait for Clk_period;
		Addr <=  "0010011100011";
		Trees_din <= x"a1ff8e04";
		wait for Clk_period;
		Addr <=  "0010011100100";
		Trees_din <= x"ffe513d9";
		wait for Clk_period;
		Addr <=  "0010011100101";
		Trees_din <= x"008613d9";
		wait for Clk_period;
		Addr <=  "0010011100110";
		Trees_din <= x"ecffb604";
		wait for Clk_period;
		Addr <=  "0010011100111";
		Trees_din <= x"004313d9";
		wait for Clk_period;
		Addr <=  "0010011101000";
		Trees_din <= x"8500a504";
		wait for Clk_period;
		Addr <=  "0010011101001";
		Trees_din <= x"ff6f13d9";
		wait for Clk_period;
		Addr <=  "0010011101010";
		Trees_din <= x"000f13d9";
		wait for Clk_period;
		Addr <=  "0010011101011";
		Trees_din <= x"eeff760c";
		wait for Clk_period;
		Addr <=  "0010011101100";
		Trees_din <= x"86ff5504";
		wait for Clk_period;
		Addr <=  "0010011101101";
		Trees_din <= x"ff9c13d9";
		wait for Clk_period;
		Addr <=  "0010011101110";
		Trees_din <= x"9cff2604";
		wait for Clk_period;
		Addr <=  "0010011101111";
		Trees_din <= x"009313d9";
		wait for Clk_period;
		Addr <=  "0010011110000";
		Trees_din <= x"001e13d9";
		wait for Clk_period;
		Addr <=  "0010011110001";
		Trees_din <= x"38fe6904";
		wait for Clk_period;
		Addr <=  "0010011110010";
		Trees_din <= x"003f13d9";
		wait for Clk_period;
		Addr <=  "0010011110011";
		Trees_din <= x"90001404";
		wait for Clk_period;
		Addr <=  "0010011110100";
		Trees_din <= x"ff6b13d9";
		wait for Clk_period;
		Addr <=  "0010011110101";
		Trees_din <= x"ffde13d9";
		wait for Clk_period;
		Addr <=  "0010011110110";
		Trees_din <= x"8dfe4b14";
		wait for Clk_period;
		Addr <=  "0010011110111";
		Trees_din <= x"d1ff6208";
		wait for Clk_period;
		Addr <=  "0010011111000";
		Trees_din <= x"4aff7e04";
		wait for Clk_period;
		Addr <=  "0010011111001";
		Trees_din <= x"ff6d149d";
		wait for Clk_period;
		Addr <=  "0010011111010";
		Trees_din <= x"ffec149d";
		wait for Clk_period;
		Addr <=  "0010011111011";
		Trees_din <= x"1fff5504";
		wait for Clk_period;
		Addr <=  "0010011111100";
		Trees_din <= x"006d149d";
		wait for Clk_period;
		Addr <=  "0010011111101";
		Trees_din <= x"f2029604";
		wait for Clk_period;
		Addr <=  "0010011111110";
		Trees_din <= x"ff9f149d";
		wait for Clk_period;
		Addr <=  "0010011111111";
		Trees_din <= x"ffec149d";
		wait for Clk_period;
		Addr <=  "0010100000000";
		Trees_din <= x"3afed020";
		wait for Clk_period;
		Addr <=  "0010100000001";
		Trees_din <= x"2a004418";
		wait for Clk_period;
		Addr <=  "0010100000010";
		Trees_din <= x"53001510";
		wait for Clk_period;
		Addr <=  "0010100000011";
		Trees_din <= x"77ff6308";
		wait for Clk_period;
		Addr <=  "0010100000100";
		Trees_din <= x"00fee404";
		wait for Clk_period;
		Addr <=  "0010100000101";
		Trees_din <= x"ffda149d";
		wait for Clk_period;
		Addr <=  "0010100000110";
		Trees_din <= x"00a0149d";
		wait for Clk_period;
		Addr <=  "0010100000111";
		Trees_din <= x"9afff804";
		wait for Clk_period;
		Addr <=  "0010100001000";
		Trees_din <= x"003b149d";
		wait for Clk_period;
		Addr <=  "0010100001001";
		Trees_din <= x"ffa0149d";
		wait for Clk_period;
		Addr <=  "0010100001010";
		Trees_din <= x"70fe6b04";
		wait for Clk_period;
		Addr <=  "0010100001011";
		Trees_din <= x"0048149d";
		wait for Clk_period;
		Addr <=  "0010100001100";
		Trees_din <= x"ff90149d";
		wait for Clk_period;
		Addr <=  "0010100001101";
		Trees_din <= x"fcffbe04";
		wait for Clk_period;
		Addr <=  "0010100001110";
		Trees_din <= x"ff85149d";
		wait for Clk_period;
		Addr <=  "0010100001111";
		Trees_din <= x"0042149d";
		wait for Clk_period;
		Addr <=  "0010100010000";
		Trees_din <= x"a1ff1c14";
		wait for Clk_period;
		Addr <=  "0010100010001";
		Trees_din <= x"6dffbd08";
		wait for Clk_period;
		Addr <=  "0010100010010";
		Trees_din <= x"83ff2204";
		wait for Clk_period;
		Addr <=  "0010100010011";
		Trees_din <= x"0099149d";
		wait for Clk_period;
		Addr <=  "0010100010100";
		Trees_din <= x"ffaa149d";
		wait for Clk_period;
		Addr <=  "0010100010101";
		Trees_din <= x"43fe8d04";
		wait for Clk_period;
		Addr <=  "0010100010110";
		Trees_din <= x"003f149d";
		wait for Clk_period;
		Addr <=  "0010100010111";
		Trees_din <= x"c8ff4e04";
		wait for Clk_period;
		Addr <=  "0010100011000";
		Trees_din <= x"0023149d";
		wait for Clk_period;
		Addr <=  "0010100011001";
		Trees_din <= x"ff6e149d";
		wait for Clk_period;
		Addr <=  "0010100011010";
		Trees_din <= x"a4ffa410";
		wait for Clk_period;
		Addr <=  "0010100011011";
		Trees_din <= x"02ff5608";
		wait for Clk_period;
		Addr <=  "0010100011100";
		Trees_din <= x"50ff7404";
		wait for Clk_period;
		Addr <=  "0010100011101";
		Trees_din <= x"ffea149d";
		wait for Clk_period;
		Addr <=  "0010100011110";
		Trees_din <= x"ff83149d";
		wait for Clk_period;
		Addr <=  "0010100011111";
		Trees_din <= x"b3ff4904";
		wait for Clk_period;
		Addr <=  "0010100100000";
		Trees_din <= x"0053149d";
		wait for Clk_period;
		Addr <=  "0010100100001";
		Trees_din <= x"ff90149d";
		wait for Clk_period;
		Addr <=  "0010100100010";
		Trees_din <= x"83ffab08";
		wait for Clk_period;
		Addr <=  "0010100100011";
		Trees_din <= x"85ff7404";
		wait for Clk_period;
		Addr <=  "0010100100100";
		Trees_din <= x"ffec149d";
		wait for Clk_period;
		Addr <=  "0010100100101";
		Trees_din <= x"005b149d";
		wait for Clk_period;
		Addr <=  "0010100100110";
		Trees_din <= x"ff8e149d";
		wait for Clk_period;
		Addr <=  "0010100100111";
		Trees_din <= x"16ff0c44";
		wait for Clk_period;
		Addr <=  "0010100101000";
		Trees_din <= x"d3fe9520";
		wait for Clk_period;
		Addr <=  "0010100101001";
		Trees_din <= x"22000d10";
		wait for Clk_period;
		Addr <=  "0010100101010";
		Trees_din <= x"d9ffca0c";
		wait for Clk_period;
		Addr <=  "0010100101011";
		Trees_din <= x"d8004904";
		wait for Clk_period;
		Addr <=  "0010100101100";
		Trees_din <= x"fff315a1";
		wait for Clk_period;
		Addr <=  "0010100101101";
		Trees_din <= x"b9fed304";
		wait for Clk_period;
		Addr <=  "0010100101110";
		Trees_din <= x"000915a1";
		wait for Clk_period;
		Addr <=  "0010100101111";
		Trees_din <= x"009d15a1";
		wait for Clk_period;
		Addr <=  "0010100110000";
		Trees_din <= x"ffb515a1";
		wait for Clk_period;
		Addr <=  "0010100110001";
		Trees_din <= x"9a004d08";
		wait for Clk_period;
		Addr <=  "0010100110010";
		Trees_din <= x"cb001e04";
		wait for Clk_period;
		Addr <=  "0010100110011";
		Trees_din <= x"ff7f15a1";
		wait for Clk_period;
		Addr <=  "0010100110100";
		Trees_din <= x"000915a1";
		wait for Clk_period;
		Addr <=  "0010100110101";
		Trees_din <= x"77fe4304";
		wait for Clk_period;
		Addr <=  "0010100110110";
		Trees_din <= x"006915a1";
		wait for Clk_period;
		Addr <=  "0010100110111";
		Trees_din <= x"000315a1";
		wait for Clk_period;
		Addr <=  "0010100111000";
		Trees_din <= x"aa001f1c";
		wait for Clk_period;
		Addr <=  "0010100111001";
		Trees_din <= x"f6fe400c";
		wait for Clk_period;
		Addr <=  "0010100111010";
		Trees_din <= x"47ff8904";
		wait for Clk_period;
		Addr <=  "0010100111011";
		Trees_din <= x"ff9f15a1";
		wait for Clk_period;
		Addr <=  "0010100111100";
		Trees_din <= x"d4ff7604";
		wait for Clk_period;
		Addr <=  "0010100111101";
		Trees_din <= x"ffdb15a1";
		wait for Clk_period;
		Addr <=  "0010100111110";
		Trees_din <= x"008015a1";
		wait for Clk_period;
		Addr <=  "0010100111111";
		Trees_din <= x"47ff1a08";
		wait for Clk_period;
		Addr <=  "0010101000000";
		Trees_din <= x"6cff0e04";
		wait for Clk_period;
		Addr <=  "0010101000001";
		Trees_din <= x"006915a1";
		wait for Clk_period;
		Addr <=  "0010101000010";
		Trees_din <= x"ffa815a1";
		wait for Clk_period;
		Addr <=  "0010101000011";
		Trees_din <= x"b3fe7b04";
		wait for Clk_period;
		Addr <=  "0010101000100";
		Trees_din <= x"000a15a1";
		wait for Clk_period;
		Addr <=  "0010101000101";
		Trees_din <= x"ff7015a1";
		wait for Clk_period;
		Addr <=  "0010101000110";
		Trees_din <= x"e4fea704";
		wait for Clk_period;
		Addr <=  "0010101000111";
		Trees_din <= x"007815a1";
		wait for Clk_period;
		Addr <=  "0010101001000";
		Trees_din <= x"ffae15a1";
		wait for Clk_period;
		Addr <=  "0010101001001";
		Trees_din <= x"b9fedb0c";
		wait for Clk_period;
		Addr <=  "0010101001010";
		Trees_din <= x"57ffcb08";
		wait for Clk_period;
		Addr <=  "0010101001011";
		Trees_din <= x"44008c04";
		wait for Clk_period;
		Addr <=  "0010101001100";
		Trees_din <= x"ff7915a1";
		wait for Clk_period;
		Addr <=  "0010101001101";
		Trees_din <= x"001215a1";
		wait for Clk_period;
		Addr <=  "0010101001110";
		Trees_din <= x"005415a1";
		wait for Clk_period;
		Addr <=  "0010101001111";
		Trees_din <= x"ecff9e14";
		wait for Clk_period;
		Addr <=  "0010101010000";
		Trees_din <= x"49ff5708";
		wait for Clk_period;
		Addr <=  "0010101010001";
		Trees_din <= x"69ff9304";
		wait for Clk_period;
		Addr <=  "0010101010010";
		Trees_din <= x"ffda15a1";
		wait for Clk_period;
		Addr <=  "0010101010011";
		Trees_din <= x"008315a1";
		wait for Clk_period;
		Addr <=  "0010101010100";
		Trees_din <= x"6bfe4504";
		wait for Clk_period;
		Addr <=  "0010101010101";
		Trees_din <= x"003c15a1";
		wait for Clk_period;
		Addr <=  "0010101010110";
		Trees_din <= x"fbff1f04";
		wait for Clk_period;
		Addr <=  "0010101010111";
		Trees_din <= x"ffdb15a1";
		wait for Clk_period;
		Addr <=  "0010101011000";
		Trees_din <= x"ff7215a1";
		wait for Clk_period;
		Addr <=  "0010101011001";
		Trees_din <= x"f8008010";
		wait for Clk_period;
		Addr <=  "0010101011010";
		Trees_din <= x"ac003408";
		wait for Clk_period;
		Addr <=  "0010101011011";
		Trees_din <= x"e5ff3f04";
		wait for Clk_period;
		Addr <=  "0010101011100";
		Trees_din <= x"006915a1";
		wait for Clk_period;
		Addr <=  "0010101011101";
		Trees_din <= x"ffb515a1";
		wait for Clk_period;
		Addr <=  "0010101011110";
		Trees_din <= x"f1ffae04";
		wait for Clk_period;
		Addr <=  "0010101011111";
		Trees_din <= x"ff8c15a1";
		wait for Clk_period;
		Addr <=  "0010101100000";
		Trees_din <= x"002315a1";
		wait for Clk_period;
		Addr <=  "0010101100001";
		Trees_din <= x"19ff9b08";
		wait for Clk_period;
		Addr <=  "0010101100010";
		Trees_din <= x"8bffc504";
		wait for Clk_period;
		Addr <=  "0010101100011";
		Trees_din <= x"003715a1";
		wait for Clk_period;
		Addr <=  "0010101100100";
		Trees_din <= x"ff8615a1";
		wait for Clk_period;
		Addr <=  "0010101100101";
		Trees_din <= x"5bff5b04";
		wait for Clk_period;
		Addr <=  "0010101100110";
		Trees_din <= x"008c15a1";
		wait for Clk_period;
		Addr <=  "0010101100111";
		Trees_din <= x"ffcf15a1";
		wait for Clk_period;
		Addr <=  "0010101101000";
		Trees_din <= x"2200b270";
		wait for Clk_period;
		Addr <=  "0010101101001";
		Trees_din <= x"6cff6438";
		wait for Clk_period;
		Addr <=  "0010101101010";
		Trees_din <= x"f6fed018";
		wait for Clk_period;
		Addr <=  "0010101101011";
		Trees_din <= x"92feca08";
		wait for Clk_period;
		Addr <=  "0010101101100";
		Trees_din <= x"cbff2204";
		wait for Clk_period;
		Addr <=  "0010101101101";
		Trees_din <= x"002116a5";
		wait for Clk_period;
		Addr <=  "0010101101110";
		Trees_din <= x"ff8e16a5";
		wait for Clk_period;
		Addr <=  "0010101101111";
		Trees_din <= x"0afffc08";
		wait for Clk_period;
		Addr <=  "0010101110000";
		Trees_din <= x"eeffb204";
		wait for Clk_period;
		Addr <=  "0010101110001";
		Trees_din <= x"005616a5";
		wait for Clk_period;
		Addr <=  "0010101110010";
		Trees_din <= x"ff8816a5";
		wait for Clk_period;
		Addr <=  "0010101110011";
		Trees_din <= x"6fffc204";
		wait for Clk_period;
		Addr <=  "0010101110100";
		Trees_din <= x"008916a5";
		wait for Clk_period;
		Addr <=  "0010101110101";
		Trees_din <= x"ffea16a5";
		wait for Clk_period;
		Addr <=  "0010101110110";
		Trees_din <= x"e3fe6910";
		wait for Clk_period;
		Addr <=  "0010101110111";
		Trees_din <= x"cbff8708";
		wait for Clk_period;
		Addr <=  "0010101111000";
		Trees_din <= x"c1fe6a04";
		wait for Clk_period;
		Addr <=  "0010101111001";
		Trees_din <= x"ffe216a5";
		wait for Clk_period;
		Addr <=  "0010101111010";
		Trees_din <= x"009816a5";
		wait for Clk_period;
		Addr <=  "0010101111011";
		Trees_din <= x"ebff0504";
		wait for Clk_period;
		Addr <=  "0010101111100";
		Trees_din <= x"ff9b16a5";
		wait for Clk_period;
		Addr <=  "0010101111101";
		Trees_din <= x"004e16a5";
		wait for Clk_period;
		Addr <=  "0010101111110";
		Trees_din <= x"8bffd108";
		wait for Clk_period;
		Addr <=  "0010101111111";
		Trees_din <= x"f0ffa604";
		wait for Clk_period;
		Addr <=  "0010110000000";
		Trees_din <= x"003916a5";
		wait for Clk_period;
		Addr <=  "0010110000001";
		Trees_din <= x"ff9e16a5";
		wait for Clk_period;
		Addr <=  "0010110000010";
		Trees_din <= x"74002c04";
		wait for Clk_period;
		Addr <=  "0010110000011";
		Trees_din <= x"ff7f16a5";
		wait for Clk_period;
		Addr <=  "0010110000100";
		Trees_din <= x"001116a5";
		wait for Clk_period;
		Addr <=  "0010110000101";
		Trees_din <= x"64ff1f20";
		wait for Clk_period;
		Addr <=  "0010110000110";
		Trees_din <= x"c5ff4b10";
		wait for Clk_period;
		Addr <=  "0010110000111";
		Trees_din <= x"81ff3e08";
		wait for Clk_period;
		Addr <=  "0010110001000";
		Trees_din <= x"50ff2804";
		wait for Clk_period;
		Addr <=  "0010110001001";
		Trees_din <= x"005e16a5";
		wait for Clk_period;
		Addr <=  "0010110001010";
		Trees_din <= x"ffcf16a5";
		wait for Clk_period;
		Addr <=  "0010110001011";
		Trees_din <= x"c8ff9604";
		wait for Clk_period;
		Addr <=  "0010110001100";
		Trees_din <= x"001a16a5";
		wait for Clk_period;
		Addr <=  "0010110001101";
		Trees_din <= x"ff7a16a5";
		wait for Clk_period;
		Addr <=  "0010110001110";
		Trees_din <= x"91fff408";
		wait for Clk_period;
		Addr <=  "0010110001111";
		Trees_din <= x"b3ff4504";
		wait for Clk_period;
		Addr <=  "0010110010000";
		Trees_din <= x"006016a5";
		wait for Clk_period;
		Addr <=  "0010110010001";
		Trees_din <= x"ff9416a5";
		wait for Clk_period;
		Addr <=  "0010110010010";
		Trees_din <= x"51000f04";
		wait for Clk_period;
		Addr <=  "0010110010011";
		Trees_din <= x"ff8416a5";
		wait for Clk_period;
		Addr <=  "0010110010100";
		Trees_din <= x"001516a5";
		wait for Clk_period;
		Addr <=  "0010110010101";
		Trees_din <= x"bd007f10";
		wait for Clk_period;
		Addr <=  "0010110010110";
		Trees_din <= x"ce002208";
		wait for Clk_period;
		Addr <=  "0010110010111";
		Trees_din <= x"2f000804";
		wait for Clk_period;
		Addr <=  "0010110011000";
		Trees_din <= x"ff6f16a5";
		wait for Clk_period;
		Addr <=  "0010110011001";
		Trees_din <= x"fffb16a5";
		wait for Clk_period;
		Addr <=  "0010110011010";
		Trees_din <= x"b8ff0304";
		wait for Clk_period;
		Addr <=  "0010110011011";
		Trees_din <= x"003516a5";
		wait for Clk_period;
		Addr <=  "0010110011100";
		Trees_din <= x"ffde16a5";
		wait for Clk_period;
		Addr <=  "0010110011101";
		Trees_din <= x"57ff9a04";
		wait for Clk_period;
		Addr <=  "0010110011110";
		Trees_din <= x"ffae16a5";
		wait for Clk_period;
		Addr <=  "0010110011111";
		Trees_din <= x"007e16a5";
		wait for Clk_period;
		Addr <=  "0010110100000";
		Trees_din <= x"75ffa20c";
		wait for Clk_period;
		Addr <=  "0010110100001";
		Trees_din <= x"8ffeef04";
		wait for Clk_period;
		Addr <=  "0010110100010";
		Trees_din <= x"ff9916a5";
		wait for Clk_period;
		Addr <=  "0010110100011";
		Trees_din <= x"adff3704";
		wait for Clk_period;
		Addr <=  "0010110100100";
		Trees_din <= x"008216a5";
		wait for Clk_period;
		Addr <=  "0010110100101";
		Trees_din <= x"000e16a5";
		wait for Clk_period;
		Addr <=  "0010110100110";
		Trees_din <= x"f2015904";
		wait for Clk_period;
		Addr <=  "0010110100111";
		Trees_din <= x"fff916a5";
		wait for Clk_period;
		Addr <=  "0010110101000";
		Trees_din <= x"ff6f16a5";
		wait for Clk_period;
		Addr <=  "0010110101001";
		Trees_din <= x"f2026c58";
		wait for Clk_period;
		Addr <=  "0010110101010";
		Trees_din <= x"41ff2c28";
		wait for Clk_period;
		Addr <=  "0010110101011";
		Trees_din <= x"81ff4f14";
		wait for Clk_period;
		Addr <=  "0010110101100";
		Trees_din <= x"65fec704";
		wait for Clk_period;
		Addr <=  "0010110101101";
		Trees_din <= x"ff991789";
		wait for Clk_period;
		Addr <=  "0010110101110";
		Trees_din <= x"b3ff3b08";
		wait for Clk_period;
		Addr <=  "0010110101111";
		Trees_din <= x"f5ff9d04";
		wait for Clk_period;
		Addr <=  "0010110110000";
		Trees_din <= x"ffaa1789";
		wait for Clk_period;
		Addr <=  "0010110110001";
		Trees_din <= x"00701789";
		wait for Clk_period;
		Addr <=  "0010110110010";
		Trees_din <= x"a6ff1904";
		wait for Clk_period;
		Addr <=  "0010110110011";
		Trees_din <= x"00281789";
		wait for Clk_period;
		Addr <=  "0010110110100";
		Trees_din <= x"ff961789";
		wait for Clk_period;
		Addr <=  "0010110110101";
		Trees_din <= x"2c009810";
		wait for Clk_period;
		Addr <=  "0010110110110";
		Trees_din <= x"35ff7408";
		wait for Clk_period;
		Addr <=  "0010110110111";
		Trees_din <= x"57002104";
		wait for Clk_period;
		Addr <=  "0010110111000";
		Trees_din <= x"ff8a1789";
		wait for Clk_period;
		Addr <=  "0010110111001";
		Trees_din <= x"00321789";
		wait for Clk_period;
		Addr <=  "0010110111010";
		Trees_din <= x"45fef804";
		wait for Clk_period;
		Addr <=  "0010110111011";
		Trees_din <= x"00551789";
		wait for Clk_period;
		Addr <=  "0010110111100";
		Trees_din <= x"ffa61789";
		wait for Clk_period;
		Addr <=  "0010110111101";
		Trees_din <= x"006d1789";
		wait for Clk_period;
		Addr <=  "0010110111110";
		Trees_din <= x"61ff8518";
		wait for Clk_period;
		Addr <=  "0010110111111";
		Trees_din <= x"47003910";
		wait for Clk_period;
		Addr <=  "0010111000000";
		Trees_din <= x"d5005808";
		wait for Clk_period;
		Addr <=  "0010111000001";
		Trees_din <= x"75007a04";
		wait for Clk_period;
		Addr <=  "0010111000010";
		Trees_din <= x"00721789";
		wait for Clk_period;
		Addr <=  "0010111000011";
		Trees_din <= x"ffb71789";
		wait for Clk_period;
		Addr <=  "0010111000100";
		Trees_din <= x"68ff9e04";
		wait for Clk_period;
		Addr <=  "0010111000101";
		Trees_din <= x"ffb61789";
		wait for Clk_period;
		Addr <=  "0010111000110";
		Trees_din <= x"00581789";
		wait for Clk_period;
		Addr <=  "0010111000111";
		Trees_din <= x"96000b04";
		wait for Clk_period;
		Addr <=  "0010111001000";
		Trees_din <= x"ff981789";
		wait for Clk_period;
		Addr <=  "0010111001001";
		Trees_din <= x"00371789";
		wait for Clk_period;
		Addr <=  "0010111001010";
		Trees_din <= x"4dfea210";
		wait for Clk_period;
		Addr <=  "0010111001011";
		Trees_din <= x"99ff2508";
		wait for Clk_period;
		Addr <=  "0010111001100";
		Trees_din <= x"deffdd04";
		wait for Clk_period;
		Addr <=  "0010111001101";
		Trees_din <= x"ffaf1789";
		wait for Clk_period;
		Addr <=  "0010111001110";
		Trees_din <= x"007a1789";
		wait for Clk_period;
		Addr <=  "0010111001111";
		Trees_din <= x"b2ff9004";
		wait for Clk_period;
		Addr <=  "0010111010000";
		Trees_din <= x"002e1789";
		wait for Clk_period;
		Addr <=  "0010111010001";
		Trees_din <= x"ff8d1789";
		wait for Clk_period;
		Addr <=  "0010111010010";
		Trees_din <= x"61001804";
		wait for Clk_period;
		Addr <=  "0010111010011";
		Trees_din <= x"ff791789";
		wait for Clk_period;
		Addr <=  "0010111010100";
		Trees_din <= x"00261789";
		wait for Clk_period;
		Addr <=  "0010111010101";
		Trees_din <= x"7afed908";
		wait for Clk_period;
		Addr <=  "0010111010110";
		Trees_din <= x"79ff5304";
		wait for Clk_period;
		Addr <=  "0010111010111";
		Trees_din <= x"ffcc1789";
		wait for Clk_period;
		Addr <=  "0010111011000";
		Trees_din <= x"007a1789";
		wait for Clk_period;
		Addr <=  "0010111011001";
		Trees_din <= x"b3fe6108";
		wait for Clk_period;
		Addr <=  "0010111011010";
		Trees_din <= x"6efff104";
		wait for Clk_period;
		Addr <=  "0010111011011";
		Trees_din <= x"00621789";
		wait for Clk_period;
		Addr <=  "0010111011100";
		Trees_din <= x"fff51789";
		wait for Clk_period;
		Addr <=  "0010111011101";
		Trees_din <= x"0eff8908";
		wait for Clk_period;
		Addr <=  "0010111011110";
		Trees_din <= x"36fea804";
		wait for Clk_period;
		Addr <=  "0010111011111";
		Trees_din <= x"00151789";
		wait for Clk_period;
		Addr <=  "0010111100000";
		Trees_din <= x"ff721789";
		wait for Clk_period;
		Addr <=  "0010111100001";
		Trees_din <= x"00241789";
		wait for Clk_period;
		Addr <=  "0010111100010";
		Trees_din <= x"d2feb62c";
		wait for Clk_period;
		Addr <=  "0010111100011";
		Trees_din <= x"dc001e14";
		wait for Clk_period;
		Addr <=  "0010111100100";
		Trees_din <= x"4ffe5e04";
		wait for Clk_period;
		Addr <=  "0010111100101";
		Trees_din <= x"00401895";
		wait for Clk_period;
		Addr <=  "0010111100110";
		Trees_din <= x"3d00bb0c";
		wait for Clk_period;
		Addr <=  "0010111100111";
		Trees_din <= x"e6007808";
		wait for Clk_period;
		Addr <=  "0010111101000";
		Trees_din <= x"63ff1304";
		wait for Clk_period;
		Addr <=  "0010111101001";
		Trees_din <= x"ffcf1895";
		wait for Clk_period;
		Addr <=  "0010111101010";
		Trees_din <= x"ff6f1895";
		wait for Clk_period;
		Addr <=  "0010111101011";
		Trees_din <= x"002b1895";
		wait for Clk_period;
		Addr <=  "0010111101100";
		Trees_din <= x"003f1895";
		wait for Clk_period;
		Addr <=  "0010111101101";
		Trees_din <= x"e9febd08";
		wait for Clk_period;
		Addr <=  "0010111101110";
		Trees_din <= x"7bffbc04";
		wait for Clk_period;
		Addr <=  "0010111101111";
		Trees_din <= x"ff8e1895";
		wait for Clk_period;
		Addr <=  "0010111110000";
		Trees_din <= x"00031895";
		wait for Clk_period;
		Addr <=  "0010111110001";
		Trees_din <= x"a1ff2804";
		wait for Clk_period;
		Addr <=  "0010111110010";
		Trees_din <= x"ffb51895";
		wait for Clk_period;
		Addr <=  "0010111110011";
		Trees_din <= x"70ff1408";
		wait for Clk_period;
		Addr <=  "0010111110100";
		Trees_din <= x"75ffe004";
		wait for Clk_period;
		Addr <=  "0010111110101";
		Trees_din <= x"00081895";
		wait for Clk_period;
		Addr <=  "0010111110110";
		Trees_din <= x"00931895";
		wait for Clk_period;
		Addr <=  "0010111110111";
		Trees_din <= x"ffd11895";
		wait for Clk_period;
		Addr <=  "0010111111000";
		Trees_din <= x"53ff7534";
		wait for Clk_period;
		Addr <=  "0010111111001";
		Trees_din <= x"afff1c14";
		wait for Clk_period;
		Addr <=  "0010111111010";
		Trees_din <= x"2dff5210";
		wait for Clk_period;
		Addr <=  "0010111111011";
		Trees_din <= x"38ff7608";
		wait for Clk_period;
		Addr <=  "0010111111100";
		Trees_din <= x"e3fe5404";
		wait for Clk_period;
		Addr <=  "0010111111101";
		Trees_din <= x"00931895";
		wait for Clk_period;
		Addr <=  "0010111111110";
		Trees_din <= x"00241895";
		wait for Clk_period;
		Addr <=  "0010111111111";
		Trees_din <= x"f700ac04";
		wait for Clk_period;
		Addr <=  "0011000000000";
		Trees_din <= x"ffac1895";
		wait for Clk_period;
		Addr <=  "0011000000001";
		Trees_din <= x"00311895";
		wait for Clk_period;
		Addr <=  "0011000000010";
		Trees_din <= x"ff951895";
		wait for Clk_period;
		Addr <=  "0011000000011";
		Trees_din <= x"14ff5110";
		wait for Clk_period;
		Addr <=  "0011000000100";
		Trees_din <= x"33ffd508";
		wait for Clk_period;
		Addr <=  "0011000000101";
		Trees_din <= x"cf00a604";
		wait for Clk_period;
		Addr <=  "0011000000110";
		Trees_din <= x"ff711895";
		wait for Clk_period;
		Addr <=  "0011000000111";
		Trees_din <= x"ffea1895";
		wait for Clk_period;
		Addr <=  "0011000001000";
		Trees_din <= x"feffb304";
		wait for Clk_period;
		Addr <=  "0011000001001";
		Trees_din <= x"ffc21895";
		wait for Clk_period;
		Addr <=  "0011000001010";
		Trees_din <= x"00451895";
		wait for Clk_period;
		Addr <=  "0011000001011";
		Trees_din <= x"40fff308";
		wait for Clk_period;
		Addr <=  "0011000001100";
		Trees_din <= x"c4ff5c04";
		wait for Clk_period;
		Addr <=  "0011000001101";
		Trees_din <= x"00701895";
		wait for Clk_period;
		Addr <=  "0011000001110";
		Trees_din <= x"ffd31895";
		wait for Clk_period;
		Addr <=  "0011000001111";
		Trees_din <= x"0a010e04";
		wait for Clk_period;
		Addr <=  "0011000010000";
		Trees_din <= x"ff9c1895";
		wait for Clk_period;
		Addr <=  "0011000010001";
		Trees_din <= x"00461895";
		wait for Clk_period;
		Addr <=  "0011000010010";
		Trees_din <= x"16fe9208";
		wait for Clk_period;
		Addr <=  "0011000010011";
		Trees_din <= x"a0ff7d04";
		wait for Clk_period;
		Addr <=  "0011000010100";
		Trees_din <= x"ff891895";
		wait for Clk_period;
		Addr <=  "0011000010101";
		Trees_din <= x"00191895";
		wait for Clk_period;
		Addr <=  "0011000010110";
		Trees_din <= x"da000110";
		wait for Clk_period;
		Addr <=  "0011000010111";
		Trees_din <= x"e4ff2a08";
		wait for Clk_period;
		Addr <=  "0011000011000";
		Trees_din <= x"15ffb804";
		wait for Clk_period;
		Addr <=  "0011000011001";
		Trees_din <= x"00691895";
		wait for Clk_period;
		Addr <=  "0011000011010";
		Trees_din <= x"00011895";
		wait for Clk_period;
		Addr <=  "0011000011011";
		Trees_din <= x"39001404";
		wait for Clk_period;
		Addr <=  "0011000011100";
		Trees_din <= x"ffa21895";
		wait for Clk_period;
		Addr <=  "0011000011101";
		Trees_din <= x"004a1895";
		wait for Clk_period;
		Addr <=  "0011000011110";
		Trees_din <= x"18ffdf08";
		wait for Clk_period;
		Addr <=  "0011000011111";
		Trees_din <= x"04001a04";
		wait for Clk_period;
		Addr <=  "0011000100000";
		Trees_din <= x"ffaa1895";
		wait for Clk_period;
		Addr <=  "0011000100001";
		Trees_din <= x"003e1895";
		wait for Clk_period;
		Addr <=  "0011000100010";
		Trees_din <= x"24ff4a04";
		wait for Clk_period;
		Addr <=  "0011000100011";
		Trees_din <= x"000d1895";
		wait for Clk_period;
		Addr <=  "0011000100100";
		Trees_din <= x"ff851895";
		wait for Clk_period;
		Addr <=  "0011000100101";
		Trees_din <= x"16ff0c3c";
		wait for Clk_period;
		Addr <=  "0011000100110";
		Trees_din <= x"d3fe9518";
		wait for Clk_period;
		Addr <=  "0011000100111";
		Trees_din <= x"5bff8814";
		wait for Clk_period;
		Addr <=  "0011000101000";
		Trees_din <= x"96ff5408";
		wait for Clk_period;
		Addr <=  "0011000101001";
		Trees_din <= x"35ffe004";
		wait for Clk_period;
		Addr <=  "0011000101010";
		Trees_din <= x"ffa11981";
		wait for Clk_period;
		Addr <=  "0011000101011";
		Trees_din <= x"00431981";
		wait for Clk_period;
		Addr <=  "0011000101100";
		Trees_din <= x"75ffe004";
		wait for Clk_period;
		Addr <=  "0011000101101";
		Trees_din <= x"ffed1981";
		wait for Clk_period;
		Addr <=  "0011000101110";
		Trees_din <= x"6cff8f04";
		wait for Clk_period;
		Addr <=  "0011000101111";
		Trees_din <= x"00841981";
		wait for Clk_period;
		Addr <=  "0011000110000";
		Trees_din <= x"00011981";
		wait for Clk_period;
		Addr <=  "0011000110001";
		Trees_din <= x"ffa81981";
		wait for Clk_period;
		Addr <=  "0011000110010";
		Trees_din <= x"aa001f1c";
		wait for Clk_period;
		Addr <=  "0011000110011";
		Trees_din <= x"57ff8a10";
		wait for Clk_period;
		Addr <=  "0011000110100";
		Trees_din <= x"b3fe6108";
		wait for Clk_period;
		Addr <=  "0011000110101";
		Trees_din <= x"ddff3b04";
		wait for Clk_period;
		Addr <=  "0011000110110";
		Trees_din <= x"ffc41981";
		wait for Clk_period;
		Addr <=  "0011000110111";
		Trees_din <= x"00561981";
		wait for Clk_period;
		Addr <=  "0011000111000";
		Trees_din <= x"96002904";
		wait for Clk_period;
		Addr <=  "0011000111001";
		Trees_din <= x"ff721981";
		wait for Clk_period;
		Addr <=  "0011000111010";
		Trees_din <= x"00201981";
		wait for Clk_period;
		Addr <=  "0011000111011";
		Trees_din <= x"3aff0608";
		wait for Clk_period;
		Addr <=  "0011000111100";
		Trees_din <= x"91ff5804";
		wait for Clk_period;
		Addr <=  "0011000111101";
		Trees_din <= x"00721981";
		wait for Clk_period;
		Addr <=  "0011000111110";
		Trees_din <= x"ffcf1981";
		wait for Clk_period;
		Addr <=  "0011000111111";
		Trees_din <= x"ffa61981";
		wait for Clk_period;
		Addr <=  "0011001000000";
		Trees_din <= x"c4fee404";
		wait for Clk_period;
		Addr <=  "0011001000001";
		Trees_din <= x"00691981";
		wait for Clk_period;
		Addr <=  "0011001000010";
		Trees_din <= x"ffde1981";
		wait for Clk_period;
		Addr <=  "0011001000011";
		Trees_din <= x"83ff3a18";
		wait for Clk_period;
		Addr <=  "0011001000100";
		Trees_din <= x"61ffda14";
		wait for Clk_period;
		Addr <=  "0011001000101";
		Trees_din <= x"e7fffb10";
		wait for Clk_period;
		Addr <=  "0011001000110";
		Trees_din <= x"bbfee508";
		wait for Clk_period;
		Addr <=  "0011001000111";
		Trees_din <= x"68ff1a04";
		wait for Clk_period;
		Addr <=  "0011001001000";
		Trees_din <= x"ff9b1981";
		wait for Clk_period;
		Addr <=  "0011001001001";
		Trees_din <= x"002f1981";
		wait for Clk_period;
		Addr <=  "0011001001010";
		Trees_din <= x"c8008004";
		wait for Clk_period;
		Addr <=  "0011001001011";
		Trees_din <= x"00531981";
		wait for Clk_period;
		Addr <=  "0011001001100";
		Trees_din <= x"ffb61981";
		wait for Clk_period;
		Addr <=  "0011001001101";
		Trees_din <= x"ff9b1981";
		wait for Clk_period;
		Addr <=  "0011001001110";
		Trees_din <= x"ff901981";
		wait for Clk_period;
		Addr <=  "0011001001111";
		Trees_din <= x"8aff5b08";
		wait for Clk_period;
		Addr <=  "0011001010000";
		Trees_din <= x"ccff5304";
		wait for Clk_period;
		Addr <=  "0011001010001";
		Trees_din <= x"fff61981";
		wait for Clk_period;
		Addr <=  "0011001010010";
		Trees_din <= x"ff841981";
		wait for Clk_period;
		Addr <=  "0011001010011";
		Trees_din <= x"14ff2e0c";
		wait for Clk_period;
		Addr <=  "0011001010100";
		Trees_din <= x"3afeba04";
		wait for Clk_period;
		Addr <=  "0011001010101";
		Trees_din <= x"00301981";
		wait for Clk_period;
		Addr <=  "0011001010110";
		Trees_din <= x"f7009704";
		wait for Clk_period;
		Addr <=  "0011001010111";
		Trees_din <= x"ff7d1981";
		wait for Clk_period;
		Addr <=  "0011001011000";
		Trees_din <= x"00161981";
		wait for Clk_period;
		Addr <=  "0011001011001";
		Trees_din <= x"37ffb408";
		wait for Clk_period;
		Addr <=  "0011001011010";
		Trees_din <= x"68fea604";
		wait for Clk_period;
		Addr <=  "0011001011011";
		Trees_din <= x"004b1981";
		wait for Clk_period;
		Addr <=  "0011001011100";
		Trees_din <= x"ffb31981";
		wait for Clk_period;
		Addr <=  "0011001011101";
		Trees_din <= x"f201f704";
		wait for Clk_period;
		Addr <=  "0011001011110";
		Trees_din <= x"00831981";
		wait for Clk_period;
		Addr <=  "0011001011111";
		Trees_din <= x"00011981";
		wait for Clk_period;
		Addr <=  "0011001100000";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0011001100001";
		Trees_din <= x"2200b24c";
		wait for Clk_period;
		Addr <=  "0011001100010";
		Trees_din <= x"2300073c";
		wait for Clk_period;
		Addr <=  "0011001100011";
		Trees_din <= x"b3ff4b20";
		wait for Clk_period;
		Addr <=  "0011001100100";
		Trees_din <= x"e0fef010";
		wait for Clk_period;
		Addr <=  "0011001100101";
		Trees_din <= x"2a003508";
		wait for Clk_period;
		Addr <=  "0011001100110";
		Trees_din <= x"e1ffeb04";
		wait for Clk_period;
		Addr <=  "0011001100111";
		Trees_din <= x"00761a39";
		wait for Clk_period;
		Addr <=  "0011001101000";
		Trees_din <= x"000c1a39";
		wait for Clk_period;
		Addr <=  "0011001101001";
		Trees_din <= x"9cff9404";
		wait for Clk_period;
		Addr <=  "0011001101010";
		Trees_din <= x"ff9e1a39";
		wait for Clk_period;
		Addr <=  "0011001101011";
		Trees_din <= x"002a1a39";
		wait for Clk_period;
		Addr <=  "0011001101100";
		Trees_din <= x"1bffd508";
		wait for Clk_period;
		Addr <=  "0011001101101";
		Trees_din <= x"53ff5d04";
		wait for Clk_period;
		Addr <=  "0011001101110";
		Trees_din <= x"ffd41a39";
		wait for Clk_period;
		Addr <=  "0011001101111";
		Trees_din <= x"00401a39";
		wait for Clk_period;
		Addr <=  "0011001110000";
		Trees_din <= x"6dffbd04";
		wait for Clk_period;
		Addr <=  "0011001110001";
		Trees_din <= x"00391a39";
		wait for Clk_period;
		Addr <=  "0011001110010";
		Trees_din <= x"ffab1a39";
		wait for Clk_period;
		Addr <=  "0011001110011";
		Trees_din <= x"63ffa10c";
		wait for Clk_period;
		Addr <=  "0011001110100";
		Trees_din <= x"edff3504";
		wait for Clk_period;
		Addr <=  "0011001110101";
		Trees_din <= x"ffff1a39";
		wait for Clk_period;
		Addr <=  "0011001110110";
		Trees_din <= x"38fed904";
		wait for Clk_period;
		Addr <=  "0011001110111";
		Trees_din <= x"fff01a39";
		wait for Clk_period;
		Addr <=  "0011001111000";
		Trees_din <= x"ff771a39";
		wait for Clk_period;
		Addr <=  "0011001111001";
		Trees_din <= x"83ff0f08";
		wait for Clk_period;
		Addr <=  "0011001111010";
		Trees_din <= x"59ffb004";
		wait for Clk_period;
		Addr <=  "0011001111011";
		Trees_din <= x"007e1a39";
		wait for Clk_period;
		Addr <=  "0011001111100";
		Trees_din <= x"fffd1a39";
		wait for Clk_period;
		Addr <=  "0011001111101";
		Trees_din <= x"beff5204";
		wait for Clk_period;
		Addr <=  "0011001111110";
		Trees_din <= x"00281a39";
		wait for Clk_period;
		Addr <=  "0011001111111";
		Trees_din <= x"ff871a39";
		wait for Clk_period;
		Addr <=  "0011010000000";
		Trees_din <= x"49fef304";
		wait for Clk_period;
		Addr <=  "0011010000001";
		Trees_din <= x"00411a39";
		wait for Clk_period;
		Addr <=  "0011010000010";
		Trees_din <= x"f6fe8c04";
		wait for Clk_period;
		Addr <=  "0011010000011";
		Trees_din <= x"fff51a39";
		wait for Clk_period;
		Addr <=  "0011010000100";
		Trees_din <= x"64ffbd04";
		wait for Clk_period;
		Addr <=  "0011010000101";
		Trees_din <= x"ff761a39";
		wait for Clk_period;
		Addr <=  "0011010000110";
		Trees_din <= x"ffe21a39";
		wait for Clk_period;
		Addr <=  "0011010000111";
		Trees_din <= x"75ffa208";
		wait for Clk_period;
		Addr <=  "0011010001000";
		Trees_din <= x"8ffeef04";
		wait for Clk_period;
		Addr <=  "0011010001001";
		Trees_din <= x"ffaa1a39";
		wait for Clk_period;
		Addr <=  "0011010001010";
		Trees_din <= x"00551a39";
		wait for Clk_period;
		Addr <=  "0011010001011";
		Trees_din <= x"beff4a04";
		wait for Clk_period;
		Addr <=  "0011010001100";
		Trees_din <= x"fff21a39";
		wait for Clk_period;
		Addr <=  "0011010001101";
		Trees_din <= x"ff751a39";
		wait for Clk_period;
		Addr <=  "0011010001110";
		Trees_din <= x"d2feb62c";
		wait for Clk_period;
		Addr <=  "0011010001111";
		Trees_din <= x"38ff1c14";
		wait for Clk_period;
		Addr <=  "0011010010000";
		Trees_din <= x"b2ffb50c";
		wait for Clk_period;
		Addr <=  "0011010010001";
		Trees_din <= x"ac001508";
		wait for Clk_period;
		Addr <=  "0011010010010";
		Trees_din <= x"44ffe404";
		wait for Clk_period;
		Addr <=  "0011010010011";
		Trees_din <= x"00801b25";
		wait for Clk_period;
		Addr <=  "0011010010100";
		Trees_din <= x"00141b25";
		wait for Clk_period;
		Addr <=  "0011010010101";
		Trees_din <= x"ffd21b25";
		wait for Clk_period;
		Addr <=  "0011010010110";
		Trees_din <= x"23fedc04";
		wait for Clk_period;
		Addr <=  "0011010010111";
		Trees_din <= x"00431b25";
		wait for Clk_period;
		Addr <=  "0011010011000";
		Trees_din <= x"ff981b25";
		wait for Clk_period;
		Addr <=  "0011010011001";
		Trees_din <= x"4dff220c";
		wait for Clk_period;
		Addr <=  "0011010011010";
		Trees_din <= x"5d005608";
		wait for Clk_period;
		Addr <=  "0011010011011";
		Trees_din <= x"f1003104";
		wait for Clk_period;
		Addr <=  "0011010011100";
		Trees_din <= x"ff701b25";
		wait for Clk_period;
		Addr <=  "0011010011101";
		Trees_din <= x"ffdc1b25";
		wait for Clk_period;
		Addr <=  "0011010011110";
		Trees_din <= x"00031b25";
		wait for Clk_period;
		Addr <=  "0011010011111";
		Trees_din <= x"83ff5c08";
		wait for Clk_period;
		Addr <=  "0011010100000";
		Trees_din <= x"4effb704";
		wait for Clk_period;
		Addr <=  "0011010100001";
		Trees_din <= x"fff01b25";
		wait for Clk_period;
		Addr <=  "0011010100010";
		Trees_din <= x"005a1b25";
		wait for Clk_period;
		Addr <=  "0011010100011";
		Trees_din <= x"ffb01b25";
		wait for Clk_period;
		Addr <=  "0011010100100";
		Trees_din <= x"49ffd118";
		wait for Clk_period;
		Addr <=  "0011010100101";
		Trees_din <= x"83ff9810";
		wait for Clk_period;
		Addr <=  "0011010100110";
		Trees_din <= x"2a00a10c";
		wait for Clk_period;
		Addr <=  "0011010100111";
		Trees_din <= x"01ff8408";
		wait for Clk_period;
		Addr <=  "0011010101000";
		Trees_din <= x"59fef804";
		wait for Clk_period;
		Addr <=  "0011010101001";
		Trees_din <= x"ffbf1b25";
		wait for Clk_period;
		Addr <=  "0011010101010";
		Trees_din <= x"00491b25";
		wait for Clk_period;
		Addr <=  "0011010101011";
		Trees_din <= x"ffa91b25";
		wait for Clk_period;
		Addr <=  "0011010101100";
		Trees_din <= x"ffa91b25";
		wait for Clk_period;
		Addr <=  "0011010101101";
		Trees_din <= x"d7006204";
		wait for Clk_period;
		Addr <=  "0011010101110";
		Trees_din <= x"ff931b25";
		wait for Clk_period;
		Addr <=  "0011010101111";
		Trees_din <= x"00041b25";
		wait for Clk_period;
		Addr <=  "0011010110000";
		Trees_din <= x"93ff7f14";
		wait for Clk_period;
		Addr <=  "0011010110001";
		Trees_din <= x"b3feaf08";
		wait for Clk_period;
		Addr <=  "0011010110010";
		Trees_din <= x"cc002204";
		wait for Clk_period;
		Addr <=  "0011010110011";
		Trees_din <= x"ffca1b25";
		wait for Clk_period;
		Addr <=  "0011010110100";
		Trees_din <= x"00711b25";
		wait for Clk_period;
		Addr <=  "0011010110101";
		Trees_din <= x"6cfe9804";
		wait for Clk_period;
		Addr <=  "0011010110110";
		Trees_din <= x"001e1b25";
		wait for Clk_period;
		Addr <=  "0011010110111";
		Trees_din <= x"b9ffd504";
		wait for Clk_period;
		Addr <=  "0011010111000";
		Trees_din <= x"ff771b25";
		wait for Clk_period;
		Addr <=  "0011010111001";
		Trees_din <= x"ffeb1b25";
		wait for Clk_period;
		Addr <=  "0011010111010";
		Trees_din <= x"8dfeec10";
		wait for Clk_period;
		Addr <=  "0011010111011";
		Trees_din <= x"0efeb508";
		wait for Clk_period;
		Addr <=  "0011010111100";
		Trees_din <= x"f1ffef04";
		wait for Clk_period;
		Addr <=  "0011010111101";
		Trees_din <= x"ff931b25";
		wait for Clk_period;
		Addr <=  "0011010111110";
		Trees_din <= x"ffff1b25";
		wait for Clk_period;
		Addr <=  "0011010111111";
		Trees_din <= x"ab006f04";
		wait for Clk_period;
		Addr <=  "0011011000000";
		Trees_din <= x"007a1b25";
		wait for Clk_period;
		Addr <=  "0011011000001";
		Trees_din <= x"ffed1b25";
		wait for Clk_period;
		Addr <=  "0011011000010";
		Trees_din <= x"6cfeed08";
		wait for Clk_period;
		Addr <=  "0011011000011";
		Trees_din <= x"41ff3f04";
		wait for Clk_period;
		Addr <=  "0011011000100";
		Trees_din <= x"ffed1b25";
		wait for Clk_period;
		Addr <=  "0011011000101";
		Trees_din <= x"005c1b25";
		wait for Clk_period;
		Addr <=  "0011011000110";
		Trees_din <= x"64fe8804";
		wait for Clk_period;
		Addr <=  "0011011000111";
		Trees_din <= x"00281b25";
		wait for Clk_period;
		Addr <=  "0011011001000";
		Trees_din <= x"ff841b25";
		wait for Clk_period;
		Addr <=  "0011011001001";
		Trees_din <= x"47004654";
		wait for Clk_period;
		Addr <=  "0011011001010";
		Trees_din <= x"18000e3c";
		wait for Clk_period;
		Addr <=  "0011011001011";
		Trees_din <= x"c4ff031c";
		wait for Clk_period;
		Addr <=  "0011011001100";
		Trees_din <= x"9fffa210";
		wait for Clk_period;
		Addr <=  "0011011001101";
		Trees_din <= x"5bffb108";
		wait for Clk_period;
		Addr <=  "0011011001110";
		Trees_din <= x"6affc804";
		wait for Clk_period;
		Addr <=  "0011011001111";
		Trees_din <= x"ffc51bf9";
		wait for Clk_period;
		Addr <=  "0011011010000";
		Trees_din <= x"00341bf9";
		wait for Clk_period;
		Addr <=  "0011011010001";
		Trees_din <= x"6cff5104";
		wait for Clk_period;
		Addr <=  "0011011010010";
		Trees_din <= x"008b1bf9";
		wait for Clk_period;
		Addr <=  "0011011010011";
		Trees_din <= x"000a1bf9";
		wait for Clk_period;
		Addr <=  "0011011010100";
		Trees_din <= x"93ff6104";
		wait for Clk_period;
		Addr <=  "0011011010101";
		Trees_din <= x"fffe1bf9";
		wait for Clk_period;
		Addr <=  "0011011010110";
		Trees_din <= x"0b004c04";
		wait for Clk_period;
		Addr <=  "0011011010111";
		Trees_din <= x"00831bf9";
		wait for Clk_period;
		Addr <=  "0011011011000";
		Trees_din <= x"000b1bf9";
		wait for Clk_period;
		Addr <=  "0011011011001";
		Trees_din <= x"63ff8810";
		wait for Clk_period;
		Addr <=  "0011011011010";
		Trees_din <= x"c1feaf08";
		wait for Clk_period;
		Addr <=  "0011011011011";
		Trees_din <= x"fcff3a04";
		wait for Clk_period;
		Addr <=  "0011011011100";
		Trees_din <= x"ffa31bf9";
		wait for Clk_period;
		Addr <=  "0011011011101";
		Trees_din <= x"00331bf9";
		wait for Clk_period;
		Addr <=  "0011011011110";
		Trees_din <= x"4ffe9c04";
		wait for Clk_period;
		Addr <=  "0011011011111";
		Trees_din <= x"fff81bf9";
		wait for Clk_period;
		Addr <=  "0011011100000";
		Trees_din <= x"ff7e1bf9";
		wait for Clk_period;
		Addr <=  "0011011100001";
		Trees_din <= x"6fff4d08";
		wait for Clk_period;
		Addr <=  "0011011100010";
		Trees_din <= x"e6ff4504";
		wait for Clk_period;
		Addr <=  "0011011100011";
		Trees_din <= x"ffbf1bf9";
		wait for Clk_period;
		Addr <=  "0011011100100";
		Trees_din <= x"005e1bf9";
		wait for Clk_period;
		Addr <=  "0011011100101";
		Trees_din <= x"e0feee04";
		wait for Clk_period;
		Addr <=  "0011011100110";
		Trees_din <= x"002e1bf9";
		wait for Clk_period;
		Addr <=  "0011011100111";
		Trees_din <= x"ffc51bf9";
		wait for Clk_period;
		Addr <=  "0011011101000";
		Trees_din <= x"02ff0308";
		wait for Clk_period;
		Addr <=  "0011011101001";
		Trees_din <= x"c6fff604";
		wait for Clk_period;
		Addr <=  "0011011101010";
		Trees_din <= x"ff791bf9";
		wait for Clk_period;
		Addr <=  "0011011101011";
		Trees_din <= x"001a1bf9";
		wait for Clk_period;
		Addr <=  "0011011101100";
		Trees_din <= x"5bff6b08";
		wait for Clk_period;
		Addr <=  "0011011101101";
		Trees_din <= x"3eff7a04";
		wait for Clk_period;
		Addr <=  "0011011101110";
		Trees_din <= x"ffa31bf9";
		wait for Clk_period;
		Addr <=  "0011011101111";
		Trees_din <= x"fffe1bf9";
		wait for Clk_period;
		Addr <=  "0011011110000";
		Trees_din <= x"eeffc504";
		wait for Clk_period;
		Addr <=  "0011011110001";
		Trees_din <= x"00641bf9";
		wait for Clk_period;
		Addr <=  "0011011110010";
		Trees_din <= x"ffef1bf9";
		wait for Clk_period;
		Addr <=  "0011011110011";
		Trees_din <= x"f1002710";
		wait for Clk_period;
		Addr <=  "0011011110100";
		Trees_din <= x"b1ff7a08";
		wait for Clk_period;
		Addr <=  "0011011110101";
		Trees_din <= x"3bfe8c04";
		wait for Clk_period;
		Addr <=  "0011011110110";
		Trees_din <= x"fffe1bf9";
		wait for Clk_period;
		Addr <=  "0011011110111";
		Trees_din <= x"ff751bf9";
		wait for Clk_period;
		Addr <=  "0011011111000";
		Trees_din <= x"7c000704";
		wait for Clk_period;
		Addr <=  "0011011111001";
		Trees_din <= x"ffd51bf9";
		wait for Clk_period;
		Addr <=  "0011011111010";
		Trees_din <= x"003f1bf9";
		wait for Clk_period;
		Addr <=  "0011011111011";
		Trees_din <= x"85000b04";
		wait for Clk_period;
		Addr <=  "0011011111100";
		Trees_din <= x"ffc31bf9";
		wait for Clk_period;
		Addr <=  "0011011111101";
		Trees_din <= x"00621bf9";
		wait for Clk_period;
		Addr <=  "0011011111110";
		Trees_din <= x"6cff6444";
		wait for Clk_period;
		Addr <=  "0011011111111";
		Trees_din <= x"6fffd138";
		wait for Clk_period;
		Addr <=  "0011100000000";
		Trees_din <= x"faff8d20";
		wait for Clk_period;
		Addr <=  "0011100000001";
		Trees_din <= x"f0ff7410";
		wait for Clk_period;
		Addr <=  "0011100000010";
		Trees_din <= x"35fea808";
		wait for Clk_period;
		Addr <=  "0011100000011";
		Trees_din <= x"15ff4704";
		wait for Clk_period;
		Addr <=  "0011100000100";
		Trees_din <= x"002a1cf5";
		wait for Clk_period;
		Addr <=  "0011100000101";
		Trees_din <= x"ffa81cf5";
		wait for Clk_period;
		Addr <=  "0011100000110";
		Trees_din <= x"efff1c04";
		wait for Clk_period;
		Addr <=  "0011100000111";
		Trees_din <= x"000b1cf5";
		wait for Clk_period;
		Addr <=  "0011100001000";
		Trees_din <= x"006b1cf5";
		wait for Clk_period;
		Addr <=  "0011100001001";
		Trees_din <= x"1eff8708";
		wait for Clk_period;
		Addr <=  "0011100001010";
		Trees_din <= x"71ff1a04";
		wait for Clk_period;
		Addr <=  "0011100001011";
		Trees_din <= x"ffe41cf5";
		wait for Clk_period;
		Addr <=  "0011100001100";
		Trees_din <= x"ff8d1cf5";
		wait for Clk_period;
		Addr <=  "0011100001101";
		Trees_din <= x"e2ff6c04";
		wait for Clk_period;
		Addr <=  "0011100001110";
		Trees_din <= x"00541cf5";
		wait for Clk_period;
		Addr <=  "0011100001111";
		Trees_din <= x"ffd51cf5";
		wait for Clk_period;
		Addr <=  "0011100010000";
		Trees_din <= x"50ff7110";
		wait for Clk_period;
		Addr <=  "0011100010001";
		Trees_din <= x"25fff608";
		wait for Clk_period;
		Addr <=  "0011100010010";
		Trees_din <= x"16ff3604";
		wait for Clk_period;
		Addr <=  "0011100010011";
		Trees_din <= x"ffe41cf5";
		wait for Clk_period;
		Addr <=  "0011100010100";
		Trees_din <= x"006d1cf5";
		wait for Clk_period;
		Addr <=  "0011100010101";
		Trees_din <= x"c9003604";
		wait for Clk_period;
		Addr <=  "0011100010110";
		Trees_din <= x"ffaf1cf5";
		wait for Clk_period;
		Addr <=  "0011100010111";
		Trees_din <= x"00311cf5";
		wait for Clk_period;
		Addr <=  "0011100011000";
		Trees_din <= x"1f002f04";
		wait for Clk_period;
		Addr <=  "0011100011001";
		Trees_din <= x"ff861cf5";
		wait for Clk_period;
		Addr <=  "0011100011010";
		Trees_din <= x"ffeb1cf5";
		wait for Clk_period;
		Addr <=  "0011100011011";
		Trees_din <= x"1cfef604";
		wait for Clk_period;
		Addr <=  "0011100011100";
		Trees_din <= x"003c1cf5";
		wait for Clk_period;
		Addr <=  "0011100011101";
		Trees_din <= x"11ffa904";
		wait for Clk_period;
		Addr <=  "0011100011110";
		Trees_din <= x"ff831cf5";
		wait for Clk_period;
		Addr <=  "0011100011111";
		Trees_din <= x"ffeb1cf5";
		wait for Clk_period;
		Addr <=  "0011100100000";
		Trees_din <= x"c5ff4b18";
		wait for Clk_period;
		Addr <=  "0011100100001";
		Trees_din <= x"3afeba0c";
		wait for Clk_period;
		Addr <=  "0011100100010";
		Trees_din <= x"d2fef804";
		wait for Clk_period;
		Addr <=  "0011100100011";
		Trees_din <= x"ffbf1cf5";
		wait for Clk_period;
		Addr <=  "0011100100100";
		Trees_din <= x"a4ffd504";
		wait for Clk_period;
		Addr <=  "0011100100101";
		Trees_din <= x"000a1cf5";
		wait for Clk_period;
		Addr <=  "0011100100110";
		Trees_din <= x"005d1cf5";
		wait for Clk_period;
		Addr <=  "0011100100111";
		Trees_din <= x"9fffb804";
		wait for Clk_period;
		Addr <=  "0011100101000";
		Trees_din <= x"ff751cf5";
		wait for Clk_period;
		Addr <=  "0011100101001";
		Trees_din <= x"0400ac04";
		wait for Clk_period;
		Addr <=  "0011100101010";
		Trees_din <= x"ffa81cf5";
		wait for Clk_period;
		Addr <=  "0011100101011";
		Trees_din <= x"004b1cf5";
		wait for Clk_period;
		Addr <=  "0011100101100";
		Trees_din <= x"9affcf0c";
		wait for Clk_period;
		Addr <=  "0011100101101";
		Trees_din <= x"abff6804";
		wait for Clk_period;
		Addr <=  "0011100101110";
		Trees_din <= x"00361cf5";
		wait for Clk_period;
		Addr <=  "0011100101111";
		Trees_din <= x"39fef404";
		wait for Clk_period;
		Addr <=  "0011100110000";
		Trees_din <= x"ffdf1cf5";
		wait for Clk_period;
		Addr <=  "0011100110001";
		Trees_din <= x"ff831cf5";
		wait for Clk_period;
		Addr <=  "0011100110010";
		Trees_din <= x"3bff6d10";
		wait for Clk_period;
		Addr <=  "0011100110011";
		Trees_din <= x"16fee708";
		wait for Clk_period;
		Addr <=  "0011100110100";
		Trees_din <= x"c3002804";
		wait for Clk_period;
		Addr <=  "0011100110101";
		Trees_din <= x"ffa01cf5";
		wait for Clk_period;
		Addr <=  "0011100110110";
		Trees_din <= x"00271cf5";
		wait for Clk_period;
		Addr <=  "0011100110111";
		Trees_din <= x"8fff6504";
		wait for Clk_period;
		Addr <=  "0011100111000";
		Trees_din <= x"00651cf5";
		wait for Clk_period;
		Addr <=  "0011100111001";
		Trees_din <= x"ffd21cf5";
		wait for Clk_period;
		Addr <=  "0011100111010";
		Trees_din <= x"1bff2f04";
		wait for Clk_period;
		Addr <=  "0011100111011";
		Trees_din <= x"002e1cf5";
		wait for Clk_period;
		Addr <=  "0011100111100";
		Trees_din <= x"ff931cf5";
		wait for Clk_period;
		Addr <=  "0011100111101";
		Trees_din <= x"47003260";
		wait for Clk_period;
		Addr <=  "0011100111110";
		Trees_din <= x"61ff8534";
		wait for Clk_period;
		Addr <=  "0011100111111";
		Trees_din <= x"63ff741c";
		wait for Clk_period;
		Addr <=  "0011101000000";
		Trees_din <= x"38ff3a10";
		wait for Clk_period;
		Addr <=  "0011101000001";
		Trees_din <= x"01feec08";
		wait for Clk_period;
		Addr <=  "0011101000010";
		Trees_din <= x"b7ffc804";
		wait for Clk_period;
		Addr <=  "0011101000011";
		Trees_din <= x"ffab1de9";
		wait for Clk_period;
		Addr <=  "0011101000100";
		Trees_din <= x"000a1de9";
		wait for Clk_period;
		Addr <=  "0011101000101";
		Trees_din <= x"22001b04";
		wait for Clk_period;
		Addr <=  "0011101000110";
		Trees_din <= x"006f1de9";
		wait for Clk_period;
		Addr <=  "0011101000111";
		Trees_din <= x"fff31de9";
		wait for Clk_period;
		Addr <=  "0011101001000";
		Trees_din <= x"b3fead04";
		wait for Clk_period;
		Addr <=  "0011101001001";
		Trees_din <= x"001b1de9";
		wait for Clk_period;
		Addr <=  "0011101001010";
		Trees_din <= x"eeff8f04";
		wait for Clk_period;
		Addr <=  "0011101001011";
		Trees_din <= x"fffc1de9";
		wait for Clk_period;
		Addr <=  "0011101001100";
		Trees_din <= x"ff831de9";
		wait for Clk_period;
		Addr <=  "0011101001101";
		Trees_din <= x"e5ff3f10";
		wait for Clk_period;
		Addr <=  "0011101001110";
		Trees_din <= x"41feb008";
		wait for Clk_period;
		Addr <=  "0011101001111";
		Trees_din <= x"61fe8f04";
		wait for Clk_period;
		Addr <=  "0011101010000";
		Trees_din <= x"00211de9";
		wait for Clk_period;
		Addr <=  "0011101010001";
		Trees_din <= x"ff9f1de9";
		wait for Clk_period;
		Addr <=  "0011101010010";
		Trees_din <= x"83ff9f04";
		wait for Clk_period;
		Addr <=  "0011101010011";
		Trees_din <= x"00561de9";
		wait for Clk_period;
		Addr <=  "0011101010100";
		Trees_din <= x"ffd71de9";
		wait for Clk_period;
		Addr <=  "0011101010101";
		Trees_din <= x"21ff6b04";
		wait for Clk_period;
		Addr <=  "0011101010110";
		Trees_din <= x"00151de9";
		wait for Clk_period;
		Addr <=  "0011101010111";
		Trees_din <= x"ff9f1de9";
		wait for Clk_period;
		Addr <=  "0011101011000";
		Trees_din <= x"97fea20c";
		wait for Clk_period;
		Addr <=  "0011101011001";
		Trees_din <= x"85000708";
		wait for Clk_period;
		Addr <=  "0011101011010";
		Trees_din <= x"55ff9304";
		wait for Clk_period;
		Addr <=  "0011101011011";
		Trees_din <= x"004e1de9";
		wait for Clk_period;
		Addr <=  "0011101011100";
		Trees_din <= x"ffb91de9";
		wait for Clk_period;
		Addr <=  "0011101011101";
		Trees_din <= x"00741de9";
		wait for Clk_period;
		Addr <=  "0011101011110";
		Trees_din <= x"27fff110";
		wait for Clk_period;
		Addr <=  "0011101011111";
		Trees_din <= x"c1fe4b08";
		wait for Clk_period;
		Addr <=  "0011101100000";
		Trees_din <= x"0cff0904";
		wait for Clk_period;
		Addr <=  "0011101100001";
		Trees_din <= x"ffcc1de9";
		wait for Clk_period;
		Addr <=  "0011101100010";
		Trees_din <= x"005b1de9";
		wait for Clk_period;
		Addr <=  "0011101100011";
		Trees_din <= x"adff2404";
		wait for Clk_period;
		Addr <=  "0011101100100";
		Trees_din <= x"fff91de9";
		wait for Clk_period;
		Addr <=  "0011101100101";
		Trees_din <= x"ff7c1de9";
		wait for Clk_period;
		Addr <=  "0011101100110";
		Trees_din <= x"05006208";
		wait for Clk_period;
		Addr <=  "0011101100111";
		Trees_din <= x"71ffbb04";
		wait for Clk_period;
		Addr <=  "0011101101000";
		Trees_din <= x"ff991de9";
		wait for Clk_period;
		Addr <=  "0011101101001";
		Trees_din <= x"00171de9";
		wait for Clk_period;
		Addr <=  "0011101101010";
		Trees_din <= x"9fff4904";
		wait for Clk_period;
		Addr <=  "0011101101011";
		Trees_din <= x"ffe41de9";
		wait for Clk_period;
		Addr <=  "0011101101100";
		Trees_din <= x"00721de9";
		wait for Clk_period;
		Addr <=  "0011101101101";
		Trees_din <= x"dcfff108";
		wait for Clk_period;
		Addr <=  "0011101101110";
		Trees_din <= x"afff1704";
		wait for Clk_period;
		Addr <=  "0011101101111";
		Trees_din <= x"fff31de9";
		wait for Clk_period;
		Addr <=  "0011101110000";
		Trees_din <= x"ff7a1de9";
		wait for Clk_period;
		Addr <=  "0011101110001";
		Trees_din <= x"d2fedc04";
		wait for Clk_period;
		Addr <=  "0011101110010";
		Trees_din <= x"ffa11de9";
		wait for Clk_period;
		Addr <=  "0011101110011";
		Trees_din <= x"7200470c";
		wait for Clk_period;
		Addr <=  "0011101110100";
		Trees_din <= x"b9ff5a08";
		wait for Clk_period;
		Addr <=  "0011101110101";
		Trees_din <= x"defff504";
		wait for Clk_period;
		Addr <=  "0011101110110";
		Trees_din <= x"00011de9";
		wait for Clk_period;
		Addr <=  "0011101110111";
		Trees_din <= x"00701de9";
		wait for Clk_period;
		Addr <=  "0011101111000";
		Trees_din <= x"ffd91de9";
		wait for Clk_period;
		Addr <=  "0011101111001";
		Trees_din <= x"ffc81de9";
		wait for Clk_period;
		Addr <=  "0011101111010";
		Trees_din <= x"2200b240";
		wait for Clk_period;
		Addr <=  "0011101111011";
		Trees_din <= x"23000730";
		wait for Clk_period;
		Addr <=  "0011101111100";
		Trees_din <= x"c4ff0318";
		wait for Clk_period;
		Addr <=  "0011101111101";
		Trees_din <= x"a6ffab10";
		wait for Clk_period;
		Addr <=  "0011101111110";
		Trees_din <= x"35fe9508";
		wait for Clk_period;
		Addr <=  "0011101111111";
		Trees_din <= x"e4fe6004";
		wait for Clk_period;
		Addr <=  "0011110000000";
		Trees_din <= x"00401e85";
		wait for Clk_period;
		Addr <=  "0011110000001";
		Trees_din <= x"ff9b1e85";
		wait for Clk_period;
		Addr <=  "0011110000010";
		Trees_din <= x"f9ff9904";
		wait for Clk_period;
		Addr <=  "0011110000011";
		Trees_din <= x"00551e85";
		wait for Clk_period;
		Addr <=  "0011110000100";
		Trees_din <= x"ffc91e85";
		wait for Clk_period;
		Addr <=  "0011110000101";
		Trees_din <= x"adff4a04";
		wait for Clk_period;
		Addr <=  "0011110000110";
		Trees_din <= x"00141e85";
		wait for Clk_period;
		Addr <=  "0011110000111";
		Trees_din <= x"ffa11e85";
		wait for Clk_period;
		Addr <=  "0011110001000";
		Trees_din <= x"53ff2a08";
		wait for Clk_period;
		Addr <=  "0011110001001";
		Trees_din <= x"8affe204";
		wait for Clk_period;
		Addr <=  "0011110001010";
		Trees_din <= x"ff8a1e85";
		wait for Clk_period;
		Addr <=  "0011110001011";
		Trees_din <= x"fff71e85";
		wait for Clk_period;
		Addr <=  "0011110001100";
		Trees_din <= x"70ff6708";
		wait for Clk_period;
		Addr <=  "0011110001101";
		Trees_din <= x"d2fecf04";
		wait for Clk_period;
		Addr <=  "0011110001110";
		Trees_din <= x"ffd81e85";
		wait for Clk_period;
		Addr <=  "0011110001111";
		Trees_din <= x"002d1e85";
		wait for Clk_period;
		Addr <=  "0011110010000";
		Trees_din <= x"9cffa704";
		wait for Clk_period;
		Addr <=  "0011110010001";
		Trees_din <= x"ff871e85";
		wait for Clk_period;
		Addr <=  "0011110010010";
		Trees_din <= x"001f1e85";
		wait for Clk_period;
		Addr <=  "0011110010011";
		Trees_din <= x"9fffda08";
		wait for Clk_period;
		Addr <=  "0011110010100";
		Trees_din <= x"34ffb104";
		wait for Clk_period;
		Addr <=  "0011110010101";
		Trees_din <= x"fff81e85";
		wait for Clk_period;
		Addr <=  "0011110010110";
		Trees_din <= x"ff7f1e85";
		wait for Clk_period;
		Addr <=  "0011110010111";
		Trees_din <= x"36ff6704";
		wait for Clk_period;
		Addr <=  "0011110011000";
		Trees_din <= x"fff01e85";
		wait for Clk_period;
		Addr <=  "0011110011001";
		Trees_din <= x"00451e85";
		wait for Clk_period;
		Addr <=  "0011110011010";
		Trees_din <= x"75ffa208";
		wait for Clk_period;
		Addr <=  "0011110011011";
		Trees_din <= x"89ffe104";
		wait for Clk_period;
		Addr <=  "0011110011100";
		Trees_din <= x"ffcd1e85";
		wait for Clk_period;
		Addr <=  "0011110011101";
		Trees_din <= x"00441e85";
		wait for Clk_period;
		Addr <=  "0011110011110";
		Trees_din <= x"93ffe104";
		wait for Clk_period;
		Addr <=  "0011110011111";
		Trees_din <= x"ff811e85";
		wait for Clk_period;
		Addr <=  "0011110100000";
		Trees_din <= x"ffdd1e85";
		wait for Clk_period;
		Addr <=  "0011110100001";
		Trees_din <= x"6cff6458";
		wait for Clk_period;
		Addr <=  "0011110100010";
		Trees_din <= x"18ffbb30";
		wait for Clk_period;
		Addr <=  "0011110100011";
		Trees_din <= x"1eff6614";
		wait for Clk_period;
		Addr <=  "0011110100100";
		Trees_din <= x"d3fe4104";
		wait for Clk_period;
		Addr <=  "0011110100101";
		Trees_din <= x"00541fa1";
		wait for Clk_period;
		Addr <=  "0011110100110";
		Trees_din <= x"d4ffa608";
		wait for Clk_period;
		Addr <=  "0011110100111";
		Trees_din <= x"49ff7804";
		wait for Clk_period;
		Addr <=  "0011110101000";
		Trees_din <= x"ffed1fa1";
		wait for Clk_period;
		Addr <=  "0011110101001";
		Trees_din <= x"ff921fa1";
		wait for Clk_period;
		Addr <=  "0011110101010";
		Trees_din <= x"91ffc904";
		wait for Clk_period;
		Addr <=  "0011110101011";
		Trees_din <= x"ffed1fa1";
		wait for Clk_period;
		Addr <=  "0011110101100";
		Trees_din <= x"003e1fa1";
		wait for Clk_period;
		Addr <=  "0011110101101";
		Trees_din <= x"28ff620c";
		wait for Clk_period;
		Addr <=  "0011110101110";
		Trees_din <= x"16feb404";
		wait for Clk_period;
		Addr <=  "0011110101111";
		Trees_din <= x"ffe91fa1";
		wait for Clk_period;
		Addr <=  "0011110110000";
		Trees_din <= x"57fec604";
		wait for Clk_period;
		Addr <=  "0011110110001";
		Trees_din <= x"fff81fa1";
		wait for Clk_period;
		Addr <=  "0011110110010";
		Trees_din <= x"006a1fa1";
		wait for Clk_period;
		Addr <=  "0011110110011";
		Trees_din <= x"80ffa808";
		wait for Clk_period;
		Addr <=  "0011110110100";
		Trees_din <= x"c7ff8904";
		wait for Clk_period;
		Addr <=  "0011110110101";
		Trees_din <= x"ff9a1fa1";
		wait for Clk_period;
		Addr <=  "0011110110110";
		Trees_din <= x"00231fa1";
		wait for Clk_period;
		Addr <=  "0011110110111";
		Trees_din <= x"bd002604";
		wait for Clk_period;
		Addr <=  "0011110111000";
		Trees_din <= x"00601fa1";
		wait for Clk_period;
		Addr <=  "0011110111001";
		Trees_din <= x"ffe41fa1";
		wait for Clk_period;
		Addr <=  "0011110111010";
		Trees_din <= x"cbff5d14";
		wait for Clk_period;
		Addr <=  "0011110111011";
		Trees_din <= x"2bffad08";
		wait for Clk_period;
		Addr <=  "0011110111100";
		Trees_din <= x"db005704";
		wait for Clk_period;
		Addr <=  "0011110111101";
		Trees_din <= x"ffad1fa1";
		wait for Clk_period;
		Addr <=  "0011110111110";
		Trees_din <= x"00151fa1";
		wait for Clk_period;
		Addr <=  "0011110111111";
		Trees_din <= x"e2ff5108";
		wait for Clk_period;
		Addr <=  "0011111000000";
		Trees_din <= x"e0ff7004";
		wait for Clk_period;
		Addr <=  "0011111000001";
		Trees_din <= x"001f1fa1";
		wait for Clk_period;
		Addr <=  "0011111000010";
		Trees_din <= x"00741fa1";
		wait for Clk_period;
		Addr <=  "0011111000011";
		Trees_din <= x"00071fa1";
		wait for Clk_period;
		Addr <=  "0011111000100";
		Trees_din <= x"3dffb70c";
		wait for Clk_period;
		Addr <=  "0011111000101";
		Trees_din <= x"89ff7e04";
		wait for Clk_period;
		Addr <=  "0011111000110";
		Trees_din <= x"ffa71fa1";
		wait for Clk_period;
		Addr <=  "0011111000111";
		Trees_din <= x"3cff0204";
		wait for Clk_period;
		Addr <=  "0011111001000";
		Trees_din <= x"ffd61fa1";
		wait for Clk_period;
		Addr <=  "0011111001001";
		Trees_din <= x"004e1fa1";
		wait for Clk_period;
		Addr <=  "0011111001010";
		Trees_din <= x"8c006204";
		wait for Clk_period;
		Addr <=  "0011111001011";
		Trees_din <= x"ff7f1fa1";
		wait for Clk_period;
		Addr <=  "0011111001100";
		Trees_din <= x"00011fa1";
		wait for Clk_period;
		Addr <=  "0011111001101";
		Trees_din <= x"64ff1f28";
		wait for Clk_period;
		Addr <=  "0011111001110";
		Trees_din <= x"b9ff3010";
		wait for Clk_period;
		Addr <=  "0011111001111";
		Trees_din <= x"84001a08";
		wait for Clk_period;
		Addr <=  "0011111010000";
		Trees_din <= x"e6fff304";
		wait for Clk_period;
		Addr <=  "0011111010001";
		Trees_din <= x"ff871fa1";
		wait for Clk_period;
		Addr <=  "0011111010010";
		Trees_din <= x"fffa1fa1";
		wait for Clk_period;
		Addr <=  "0011111010011";
		Trees_din <= x"a0ff5404";
		wait for Clk_period;
		Addr <=  "0011111010100";
		Trees_din <= x"ffd41fa1";
		wait for Clk_period;
		Addr <=  "0011111010101";
		Trees_din <= x"003d1fa1";
		wait for Clk_period;
		Addr <=  "0011111010110";
		Trees_din <= x"cdffe910";
		wait for Clk_period;
		Addr <=  "0011111010111";
		Trees_din <= x"c5ff4b08";
		wait for Clk_period;
		Addr <=  "0011111011000";
		Trees_din <= x"50ff2804";
		wait for Clk_period;
		Addr <=  "0011111011001";
		Trees_din <= x"00371fa1";
		wait for Clk_period;
		Addr <=  "0011111011010";
		Trees_din <= x"ffa91fa1";
		wait for Clk_period;
		Addr <=  "0011111011011";
		Trees_din <= x"db003a04";
		wait for Clk_period;
		Addr <=  "0011111011100";
		Trees_din <= x"00711fa1";
		wait for Clk_period;
		Addr <=  "0011111011101";
		Trees_din <= x"fff11fa1";
		wait for Clk_period;
		Addr <=  "0011111011110";
		Trees_din <= x"17ffd704";
		wait for Clk_period;
		Addr <=  "0011111011111";
		Trees_din <= x"00241fa1";
		wait for Clk_period;
		Addr <=  "0011111100000";
		Trees_din <= x"ff941fa1";
		wait for Clk_period;
		Addr <=  "0011111100001";
		Trees_din <= x"beff6204";
		wait for Clk_period;
		Addr <=  "0011111100010";
		Trees_din <= x"00111fa1";
		wait for Clk_period;
		Addr <=  "0011111100011";
		Trees_din <= x"edff5908";
		wait for Clk_period;
		Addr <=  "0011111100100";
		Trees_din <= x"c2ff2e04";
		wait for Clk_period;
		Addr <=  "0011111100101";
		Trees_din <= x"00261fa1";
		wait for Clk_period;
		Addr <=  "0011111100110";
		Trees_din <= x"ffb71fa1";
		wait for Clk_period;
		Addr <=  "0011111100111";
		Trees_din <= x"ff7d1fa1";
		wait for Clk_period;
		Addr <=  "0011111101000";
		Trees_din <= x"41ff2140";
		wait for Clk_period;
		Addr <=  "0011111101001";
		Trees_din <= x"fbffc428";
		wait for Clk_period;
		Addr <=  "0011111101010";
		Trees_din <= x"8e004d20";
		wait for Clk_period;
		Addr <=  "0011111101011";
		Trees_din <= x"f6fed810";
		wait for Clk_period;
		Addr <=  "0011111101100";
		Trees_din <= x"68fec608";
		wait for Clk_period;
		Addr <=  "0011111101101";
		Trees_din <= x"68fe5404";
		wait for Clk_period;
		Addr <=  "0011111101110";
		Trees_din <= x"0000207d";
		wait for Clk_period;
		Addr <=  "0011111101111";
		Trees_din <= x"0075207d";
		wait for Clk_period;
		Addr <=  "0011111110000";
		Trees_din <= x"beff0904";
		wait for Clk_period;
		Addr <=  "0011111110001";
		Trees_din <= x"0051207d";
		wait for Clk_period;
		Addr <=  "0011111110010";
		Trees_din <= x"ffbc207d";
		wait for Clk_period;
		Addr <=  "0011111110011";
		Trees_din <= x"d7007408";
		wait for Clk_period;
		Addr <=  "0011111110100";
		Trees_din <= x"7bffc204";
		wait for Clk_period;
		Addr <=  "0011111110101";
		Trees_din <= x"ff8c207d";
		wait for Clk_period;
		Addr <=  "0011111110110";
		Trees_din <= x"001d207d";
		wait for Clk_period;
		Addr <=  "0011111110111";
		Trees_din <= x"50ff4904";
		wait for Clk_period;
		Addr <=  "0011111111000";
		Trees_din <= x"0047207d";
		wait for Clk_period;
		Addr <=  "0011111111001";
		Trees_din <= x"ffcf207d";
		wait for Clk_period;
		Addr <=  "0011111111010";
		Trees_din <= x"99ff4304";
		wait for Clk_period;
		Addr <=  "0011111111011";
		Trees_din <= x"ff95207d";
		wait for Clk_period;
		Addr <=  "0011111111100";
		Trees_din <= x"ffea207d";
		wait for Clk_period;
		Addr <=  "0011111111101";
		Trees_din <= x"45fe8408";
		wait for Clk_period;
		Addr <=  "0011111111110";
		Trees_din <= x"8effc704";
		wait for Clk_period;
		Addr <=  "0011111111111";
		Trees_din <= x"004b207d";
		wait for Clk_period;
		Addr <=  "0100000000000";
		Trees_din <= x"ffe4207d";
		wait for Clk_period;
		Addr <=  "0100000000001";
		Trees_din <= x"02ff3c08";
		wait for Clk_period;
		Addr <=  "0100000000010";
		Trees_din <= x"f700c704";
		wait for Clk_period;
		Addr <=  "0100000000011";
		Trees_din <= x"ff7e207d";
		wait for Clk_period;
		Addr <=  "0100000000100";
		Trees_din <= x"ffe4207d";
		wait for Clk_period;
		Addr <=  "0100000000101";
		Trees_din <= x"c4ff0304";
		wait for Clk_period;
		Addr <=  "0100000000110";
		Trees_din <= x"003a207d";
		wait for Clk_period;
		Addr <=  "0100000000111";
		Trees_din <= x"ffb4207d";
		wait for Clk_period;
		Addr <=  "0100000001000";
		Trees_din <= x"f9ff6b20";
		wait for Clk_period;
		Addr <=  "0100000001001";
		Trees_din <= x"01fe8b08";
		wait for Clk_period;
		Addr <=  "0100000001010";
		Trees_din <= x"a1ff8804";
		wait for Clk_period;
		Addr <=  "0100000001011";
		Trees_din <= x"ff9a207d";
		wait for Clk_period;
		Addr <=  "0100000001100";
		Trees_din <= x"001b207d";
		wait for Clk_period;
		Addr <=  "0100000001101";
		Trees_din <= x"c4ffa110";
		wait for Clk_period;
		Addr <=  "0100000001110";
		Trees_din <= x"8ffe9f08";
		wait for Clk_period;
		Addr <=  "0100000001111";
		Trees_din <= x"ebff4204";
		wait for Clk_period;
		Addr <=  "0100000010000";
		Trees_din <= x"ffac207d";
		wait for Clk_period;
		Addr <=  "0100000010001";
		Trees_din <= x"0036207d";
		wait for Clk_period;
		Addr <=  "0100000010010";
		Trees_din <= x"2c003b04";
		wait for Clk_period;
		Addr <=  "0100000010011";
		Trees_din <= x"0058207d";
		wait for Clk_period;
		Addr <=  "0100000010100";
		Trees_din <= x"ffdb207d";
		wait for Clk_period;
		Addr <=  "0100000010101";
		Trees_din <= x"2cff8b04";
		wait for Clk_period;
		Addr <=  "0100000010110";
		Trees_din <= x"001a207d";
		wait for Clk_period;
		Addr <=  "0100000010111";
		Trees_din <= x"ffa4207d";
		wait for Clk_period;
		Addr <=  "0100000011000";
		Trees_din <= x"20ff2308";
		wait for Clk_period;
		Addr <=  "0100000011001";
		Trees_din <= x"9fff9104";
		wait for Clk_period;
		Addr <=  "0100000011010";
		Trees_din <= x"fffd207d";
		wait for Clk_period;
		Addr <=  "0100000011011";
		Trees_din <= x"004b207d";
		wait for Clk_period;
		Addr <=  "0100000011100";
		Trees_din <= x"04007004";
		wait for Clk_period;
		Addr <=  "0100000011101";
		Trees_din <= x"ff8c207d";
		wait for Clk_period;
		Addr <=  "0100000011110";
		Trees_din <= x"fff1207d";
		wait for Clk_period;
		Addr <=  "0100000011111";
		Trees_din <= x"16feb214";
		wait for Clk_period;
		Addr <=  "0100000100000";
		Trees_din <= x"a0ff5408";
		wait for Clk_period;
		Addr <=  "0100000100001";
		Trees_din <= x"0bff4904";
		wait for Clk_period;
		Addr <=  "0100000100010";
		Trees_din <= x"fffc2109";
		wait for Clk_period;
		Addr <=  "0100000100011";
		Trees_din <= x"ff812109";
		wait for Clk_period;
		Addr <=  "0100000100100";
		Trees_din <= x"7aff6508";
		wait for Clk_period;
		Addr <=  "0100000100101";
		Trees_din <= x"d3fe8e04";
		wait for Clk_period;
		Addr <=  "0100000100110";
		Trees_din <= x"004e2109";
		wait for Clk_period;
		Addr <=  "0100000100111";
		Trees_din <= x"00062109";
		wait for Clk_period;
		Addr <=  "0100000101000";
		Trees_din <= x"ffc22109";
		wait for Clk_period;
		Addr <=  "0100000101001";
		Trees_din <= x"ecff9814";
		wait for Clk_period;
		Addr <=  "0100000101010";
		Trees_din <= x"c1fe7a08";
		wait for Clk_period;
		Addr <=  "0100000101011";
		Trees_din <= x"1fffb704";
		wait for Clk_period;
		Addr <=  "0100000101100";
		Trees_din <= x"ffdf2109";
		wait for Clk_period;
		Addr <=  "0100000101101";
		Trees_din <= x"004a2109";
		wait for Clk_period;
		Addr <=  "0100000101110";
		Trees_din <= x"0a00a304";
		wait for Clk_period;
		Addr <=  "0100000101111";
		Trees_din <= x"ff8a2109";
		wait for Clk_period;
		Addr <=  "0100000110000";
		Trees_din <= x"09ffd704";
		wait for Clk_period;
		Addr <=  "0100000110001";
		Trees_din <= x"ffe12109";
		wait for Clk_period;
		Addr <=  "0100000110010";
		Trees_din <= x"00262109";
		wait for Clk_period;
		Addr <=  "0100000110011";
		Trees_din <= x"c4ffd118";
		wait for Clk_period;
		Addr <=  "0100000110100";
		Trees_din <= x"6fffec10";
		wait for Clk_period;
		Addr <=  "0100000110101";
		Trees_din <= x"19ff2408";
		wait for Clk_period;
		Addr <=  "0100000110110";
		Trees_din <= x"acfff904";
		wait for Clk_period;
		Addr <=  "0100000110111";
		Trees_din <= x"00282109";
		wait for Clk_period;
		Addr <=  "0100000111000";
		Trees_din <= x"ffb02109";
		wait for Clk_period;
		Addr <=  "0100000111001";
		Trees_din <= x"cbffce04";
		wait for Clk_period;
		Addr <=  "0100000111010";
		Trees_din <= x"00402109";
		wait for Clk_period;
		Addr <=  "0100000111011";
		Trees_din <= x"fffb2109";
		wait for Clk_period;
		Addr <=  "0100000111100";
		Trees_din <= x"63ffc304";
		wait for Clk_period;
		Addr <=  "0100000111101";
		Trees_din <= x"ff972109";
		wait for Clk_period;
		Addr <=  "0100000111110";
		Trees_din <= x"000d2109";
		wait for Clk_period;
		Addr <=  "0100000111111";
		Trees_din <= x"24ffea04";
		wait for Clk_period;
		Addr <=  "0100001000000";
		Trees_din <= x"ff9c2109";
		wait for Clk_period;
		Addr <=  "0100001000001";
		Trees_din <= x"ffe82109";
		wait for Clk_period;
		Addr <=  "0100001000010";
		Trees_din <= x"41ff2134";
		wait for Clk_period;
		Addr <=  "0100001000011";
		Trees_din <= x"fbffc41c";
		wait for Clk_period;
		Addr <=  "0100001000100";
		Trees_din <= x"8e004d14";
		wait for Clk_period;
		Addr <=  "0100001000101";
		Trees_din <= x"5efff90c";
		wait for Clk_period;
		Addr <=  "0100001000110";
		Trees_din <= x"d4ff0604";
		wait for Clk_period;
		Addr <=  "0100001000111";
		Trees_din <= x"ffb621cd";
		wait for Clk_period;
		Addr <=  "0100001001000";
		Trees_din <= x"54ffef04";
		wait for Clk_period;
		Addr <=  "0100001001001";
		Trees_din <= x"ffe721cd";
		wait for Clk_period;
		Addr <=  "0100001001010";
		Trees_din <= x"004821cd";
		wait for Clk_period;
		Addr <=  "0100001001011";
		Trees_din <= x"e9fe6904";
		wait for Clk_period;
		Addr <=  "0100001001100";
		Trees_din <= x"002721cd";
		wait for Clk_period;
		Addr <=  "0100001001101";
		Trees_din <= x"ffa321cd";
		wait for Clk_period;
		Addr <=  "0100001001110";
		Trees_din <= x"6bfe7204";
		wait for Clk_period;
		Addr <=  "0100001001111";
		Trees_din <= x"fff121cd";
		wait for Clk_period;
		Addr <=  "0100001010000";
		Trees_din <= x"ff9721cd";
		wait for Clk_period;
		Addr <=  "0100001010001";
		Trees_din <= x"45fe8408";
		wait for Clk_period;
		Addr <=  "0100001010010";
		Trees_din <= x"cafe8d04";
		wait for Clk_period;
		Addr <=  "0100001010011";
		Trees_din <= x"fff921cd";
		wait for Clk_period;
		Addr <=  "0100001010100";
		Trees_din <= x"002b21cd";
		wait for Clk_period;
		Addr <=  "0100001010101";
		Trees_din <= x"5bffb90c";
		wait for Clk_period;
		Addr <=  "0100001010110";
		Trees_din <= x"a3ff0204";
		wait for Clk_period;
		Addr <=  "0100001010111";
		Trees_din <= x"ffed21cd";
		wait for Clk_period;
		Addr <=  "0100001011000";
		Trees_din <= x"f6fe4004";
		wait for Clk_period;
		Addr <=  "0100001011001";
		Trees_din <= x"ffdf21cd";
		wait for Clk_period;
		Addr <=  "0100001011010";
		Trees_din <= x"ff7b21cd";
		wait for Clk_period;
		Addr <=  "0100001011011";
		Trees_din <= x"000421cd";
		wait for Clk_period;
		Addr <=  "0100001011100";
		Trees_din <= x"18000e28";
		wait for Clk_period;
		Addr <=  "0100001011101";
		Trees_din <= x"4700251c";
		wait for Clk_period;
		Addr <=  "0100001011110";
		Trees_din <= x"f0ff6b0c";
		wait for Clk_period;
		Addr <=  "0100001011111";
		Trees_din <= x"65ffc008";
		wait for Clk_period;
		Addr <=  "0100001100000";
		Trees_din <= x"c4ff9504";
		wait for Clk_period;
		Addr <=  "0100001100001";
		Trees_din <= x"006621cd";
		wait for Clk_period;
		Addr <=  "0100001100010";
		Trees_din <= x"fff921cd";
		wait for Clk_period;
		Addr <=  "0100001100011";
		Trees_din <= x"ffe821cd";
		wait for Clk_period;
		Addr <=  "0100001100100";
		Trees_din <= x"60ff4608";
		wait for Clk_period;
		Addr <=  "0100001100101";
		Trees_din <= x"07006a04";
		wait for Clk_period;
		Addr <=  "0100001100110";
		Trees_din <= x"ff9521cd";
		wait for Clk_period;
		Addr <=  "0100001100111";
		Trees_din <= x"001b21cd";
		wait for Clk_period;
		Addr <=  "0100001101000";
		Trees_din <= x"a1ff3504";
		wait for Clk_period;
		Addr <=  "0100001101001";
		Trees_din <= x"ffbc21cd";
		wait for Clk_period;
		Addr <=  "0100001101010";
		Trees_din <= x"003621cd";
		wait for Clk_period;
		Addr <=  "0100001101011";
		Trees_din <= x"f1002708";
		wait for Clk_period;
		Addr <=  "0100001101100";
		Trees_din <= x"05000904";
		wait for Clk_period;
		Addr <=  "0100001101101";
		Trees_din <= x"000221cd";
		wait for Clk_period;
		Addr <=  "0100001101110";
		Trees_din <= x"ff9021cd";
		wait for Clk_period;
		Addr <=  "0100001101111";
		Trees_din <= x"003821cd";
		wait for Clk_period;
		Addr <=  "0100001110000";
		Trees_din <= x"34ffc304";
		wait for Clk_period;
		Addr <=  "0100001110001";
		Trees_din <= x"002021cd";
		wait for Clk_period;
		Addr <=  "0100001110010";
		Trees_din <= x"ff9b21cd";
		wait for Clk_period;
		Addr <=  "0100001110011";
		Trees_din <= x"f2026c4c";
		wait for Clk_period;
		Addr <=  "0100001110100";
		Trees_din <= x"f0ff9a30";
		wait for Clk_period;
		Addr <=  "0100001110101";
		Trees_din <= x"faff8d18";
		wait for Clk_period;
		Addr <=  "0100001110110";
		Trees_din <= x"16feb208";
		wait for Clk_period;
		Addr <=  "0100001110111";
		Trees_din <= x"5bff2404";
		wait for Clk_period;
		Addr <=  "0100001111000";
		Trees_din <= x"00212289";
		wait for Clk_period;
		Addr <=  "0100001111001";
		Trees_din <= x"ffae2289";
		wait for Clk_period;
		Addr <=  "0100001111010";
		Trees_din <= x"89ffa208";
		wait for Clk_period;
		Addr <=  "0100001111011";
		Trees_din <= x"3aff1804";
		wait for Clk_period;
		Addr <=  "0100001111100";
		Trees_din <= x"00462289";
		wait for Clk_period;
		Addr <=  "0100001111101";
		Trees_din <= x"ffcd2289";
		wait for Clk_period;
		Addr <=  "0100001111110";
		Trees_din <= x"bbff0304";
		wait for Clk_period;
		Addr <=  "0100001111111";
		Trees_din <= x"ffef2289";
		wait for Clk_period;
		Addr <=  "0100010000000";
		Trees_din <= x"00512289";
		wait for Clk_period;
		Addr <=  "0100010000001";
		Trees_din <= x"50fed708";
		wait for Clk_period;
		Addr <=  "0100010000010";
		Trees_din <= x"e8ff7904";
		wait for Clk_period;
		Addr <=  "0100010000011";
		Trees_din <= x"004d2289";
		wait for Clk_period;
		Addr <=  "0100010000100";
		Trees_din <= x"000f2289";
		wait for Clk_period;
		Addr <=  "0100010000101";
		Trees_din <= x"a9ff2708";
		wait for Clk_period;
		Addr <=  "0100010000110";
		Trees_din <= x"80ff4b04";
		wait for Clk_period;
		Addr <=  "0100010000111";
		Trees_din <= x"004e2289";
		wait for Clk_period;
		Addr <=  "0100010001000";
		Trees_din <= x"fff52289";
		wait for Clk_period;
		Addr <=  "0100010001001";
		Trees_din <= x"57001204";
		wait for Clk_period;
		Addr <=  "0100010001010";
		Trees_din <= x"ff962289";
		wait for Clk_period;
		Addr <=  "0100010001011";
		Trees_din <= x"001d2289";
		wait for Clk_period;
		Addr <=  "0100010001100";
		Trees_din <= x"2dfec00c";
		wait for Clk_period;
		Addr <=  "0100010001101";
		Trees_din <= x"b9ff6604";
		wait for Clk_period;
		Addr <=  "0100010001110";
		Trees_din <= x"ffc42289";
		wait for Clk_period;
		Addr <=  "0100010001111";
		Trees_din <= x"9a001504";
		wait for Clk_period;
		Addr <=  "0100010010000";
		Trees_din <= x"fffb2289";
		wait for Clk_period;
		Addr <=  "0100010010001";
		Trees_din <= x"005f2289";
		wait for Clk_period;
		Addr <=  "0100010010010";
		Trees_din <= x"96001d0c";
		wait for Clk_period;
		Addr <=  "0100010010011";
		Trees_din <= x"3afec204";
		wait for Clk_period;
		Addr <=  "0100010010100";
		Trees_din <= x"fffe2289";
		wait for Clk_period;
		Addr <=  "0100010010101";
		Trees_din <= x"53ff1204";
		wait for Clk_period;
		Addr <=  "0100010010110";
		Trees_din <= x"ffe72289";
		wait for Clk_period;
		Addr <=  "0100010010111";
		Trees_din <= x"ff802289";
		wait for Clk_period;
		Addr <=  "0100010011000";
		Trees_din <= x"00242289";
		wait for Clk_period;
		Addr <=  "0100010011001";
		Trees_din <= x"98fe8b0c";
		wait for Clk_period;
		Addr <=  "0100010011010";
		Trees_din <= x"d5ffd208";
		wait for Clk_period;
		Addr <=  "0100010011011";
		Trees_din <= x"c8ffe104";
		wait for Clk_period;
		Addr <=  "0100010011100";
		Trees_din <= x"00532289";
		wait for Clk_period;
		Addr <=  "0100010011101";
		Trees_din <= x"fff12289";
		wait for Clk_period;
		Addr <=  "0100010011110";
		Trees_din <= x"ffb42289";
		wait for Clk_period;
		Addr <=  "0100010011111";
		Trees_din <= x"f4ff6404";
		wait for Clk_period;
		Addr <=  "0100010100000";
		Trees_din <= x"ff872289";
		wait for Clk_period;
		Addr <=  "0100010100001";
		Trees_din <= x"000d2289";
		wait for Clk_period;
		Addr <=  "0100010100010";
		Trees_din <= x"16ff1330";
		wait for Clk_period;
		Addr <=  "0100010100011";
		Trees_din <= x"d3fe9514";
		wait for Clk_period;
		Addr <=  "0100010100100";
		Trees_din <= x"5bff8810";
		wait for Clk_period;
		Addr <=  "0100010100101";
		Trees_din <= x"f8001e04";
		wait for Clk_period;
		Addr <=  "0100010100110";
		Trees_din <= x"ffe42345";
		wait for Clk_period;
		Addr <=  "0100010100111";
		Trees_din <= x"51ffae04";
		wait for Clk_period;
		Addr <=  "0100010101000";
		Trees_din <= x"00032345";
		wait for Clk_period;
		Addr <=  "0100010101001";
		Trees_din <= x"3dfffa04";
		wait for Clk_period;
		Addr <=  "0100010101010";
		Trees_din <= x"001c2345";
		wait for Clk_period;
		Addr <=  "0100010101011";
		Trees_din <= x"00672345";
		wait for Clk_period;
		Addr <=  "0100010101100";
		Trees_din <= x"ffc52345";
		wait for Clk_period;
		Addr <=  "0100010101101";
		Trees_din <= x"23ff480c";
		wait for Clk_period;
		Addr <=  "0100010101110";
		Trees_din <= x"00ff5404";
		wait for Clk_period;
		Addr <=  "0100010101111";
		Trees_din <= x"ffb02345";
		wait for Clk_period;
		Addr <=  "0100010110000";
		Trees_din <= x"cbff9604";
		wait for Clk_period;
		Addr <=  "0100010110001";
		Trees_din <= x"00522345";
		wait for Clk_period;
		Addr <=  "0100010110010";
		Trees_din <= x"fff42345";
		wait for Clk_period;
		Addr <=  "0100010110011";
		Trees_din <= x"adff4208";
		wait for Clk_period;
		Addr <=  "0100010110100";
		Trees_din <= x"2bff6a04";
		wait for Clk_period;
		Addr <=  "0100010110101";
		Trees_din <= x"00262345";
		wait for Clk_period;
		Addr <=  "0100010110110";
		Trees_din <= x"ffc12345";
		wait for Clk_period;
		Addr <=  "0100010110111";
		Trees_din <= x"3dff7d04";
		wait for Clk_period;
		Addr <=  "0100010111000";
		Trees_din <= x"ffe52345";
		wait for Clk_period;
		Addr <=  "0100010111001";
		Trees_din <= x"ff842345";
		wait for Clk_period;
		Addr <=  "0100010111010";
		Trees_din <= x"3bffb72c";
		wait for Clk_period;
		Addr <=  "0100010111011";
		Trees_din <= x"ecff9e0c";
		wait for Clk_period;
		Addr <=  "0100010111100";
		Trees_din <= x"16ff8104";
		wait for Clk_period;
		Addr <=  "0100010111101";
		Trees_din <= x"ff9d2345";
		wait for Clk_period;
		Addr <=  "0100010111110";
		Trees_din <= x"d5ffcd04";
		wait for Clk_period;
		Addr <=  "0100010111111";
		Trees_din <= x"004c2345";
		wait for Clk_period;
		Addr <=  "0100011000000";
		Trees_din <= x"ffe82345";
		wait for Clk_period;
		Addr <=  "0100011000001";
		Trees_din <= x"f8008010";
		wait for Clk_period;
		Addr <=  "0100011000010";
		Trees_din <= x"5bff7b08";
		wait for Clk_period;
		Addr <=  "0100011000011";
		Trees_din <= x"57ffe004";
		wait for Clk_period;
		Addr <=  "0100011000100";
		Trees_din <= x"00032345";
		wait for Clk_period;
		Addr <=  "0100011000101";
		Trees_din <= x"005f2345";
		wait for Clk_period;
		Addr <=  "0100011000110";
		Trees_din <= x"20ffd504";
		wait for Clk_period;
		Addr <=  "0100011000111";
		Trees_din <= x"006a2345";
		wait for Clk_period;
		Addr <=  "0100011001000";
		Trees_din <= x"00002345";
		wait for Clk_period;
		Addr <=  "0100011001001";
		Trees_din <= x"b6ff9e08";
		wait for Clk_period;
		Addr <=  "0100011001010";
		Trees_din <= x"8bffc104";
		wait for Clk_period;
		Addr <=  "0100011001011";
		Trees_din <= x"00132345";
		wait for Clk_period;
		Addr <=  "0100011001100";
		Trees_din <= x"ffa02345";
		wait for Clk_period;
		Addr <=  "0100011001101";
		Trees_din <= x"2eff9204";
		wait for Clk_period;
		Addr <=  "0100011001110";
		Trees_din <= x"004a2345";
		wait for Clk_period;
		Addr <=  "0100011001111";
		Trees_din <= x"fff42345";
		wait for Clk_period;
		Addr <=  "0100011010000";
		Trees_din <= x"ffad2345";
		wait for Clk_period;
		Addr <=  "0100011010001";
		Trees_din <= x"f700d63c";
		wait for Clk_period;
		Addr <=  "0100011010010";
		Trees_din <= x"7affd82c";
		wait for Clk_period;
		Addr <=  "0100011010011";
		Trees_din <= x"81ff4f10";
		wait for Clk_period;
		Addr <=  "0100011010100";
		Trees_din <= x"7cffee0c";
		wait for Clk_period;
		Addr <=  "0100011010101";
		Trees_din <= x"cafdc904";
		wait for Clk_period;
		Addr <=  "0100011010110";
		Trees_din <= x"ffc923d9";
		wait for Clk_period;
		Addr <=  "0100011010111";
		Trees_din <= x"4bff2a04";
		wait for Clk_period;
		Addr <=  "0100011011000";
		Trees_din <= x"005723d9";
		wait for Clk_period;
		Addr <=  "0100011011001";
		Trees_din <= x"fff223d9";
		wait for Clk_period;
		Addr <=  "0100011011010";
		Trees_din <= x"ffbb23d9";
		wait for Clk_period;
		Addr <=  "0100011011011";
		Trees_din <= x"61ff0c0c";
		wait for Clk_period;
		Addr <=  "0100011011100";
		Trees_din <= x"c7ff0204";
		wait for Clk_period;
		Addr <=  "0100011011101";
		Trees_din <= x"ffcc23d9";
		wait for Clk_period;
		Addr <=  "0100011011110";
		Trees_din <= x"a0fee404";
		wait for Clk_period;
		Addr <=  "0100011011111";
		Trees_din <= x"ffe823d9";
		wait for Clk_period;
		Addr <=  "0100011100000";
		Trees_din <= x"004a23d9";
		wait for Clk_period;
		Addr <=  "0100011100001";
		Trees_din <= x"afff6908";
		wait for Clk_period;
		Addr <=  "0100011100010";
		Trees_din <= x"14fefd04";
		wait for Clk_period;
		Addr <=  "0100011100011";
		Trees_din <= x"ffc223d9";
		wait for Clk_period;
		Addr <=  "0100011100100";
		Trees_din <= x"003a23d9";
		wait for Clk_period;
		Addr <=  "0100011100101";
		Trees_din <= x"5ffee304";
		wait for Clk_period;
		Addr <=  "0100011100110";
		Trees_din <= x"000823d9";
		wait for Clk_period;
		Addr <=  "0100011100111";
		Trees_din <= x"ffa323d9";
		wait for Clk_period;
		Addr <=  "0100011101000";
		Trees_din <= x"d2ff4008";
		wait for Clk_period;
		Addr <=  "0100011101001";
		Trees_din <= x"ed000604";
		wait for Clk_period;
		Addr <=  "0100011101010";
		Trees_din <= x"ff8323d9";
		wait for Clk_period;
		Addr <=  "0100011101011";
		Trees_din <= x"ffdb23d9";
		wait for Clk_period;
		Addr <=  "0100011101100";
		Trees_din <= x"09febd04";
		wait for Clk_period;
		Addr <=  "0100011101101";
		Trees_din <= x"004623d9";
		wait for Clk_period;
		Addr <=  "0100011101110";
		Trees_din <= x"ffd523d9";
		wait for Clk_period;
		Addr <=  "0100011101111";
		Trees_din <= x"e3fe640c";
		wait for Clk_period;
		Addr <=  "0100011110000";
		Trees_din <= x"15ff9c04";
		wait for Clk_period;
		Addr <=  "0100011110001";
		Trees_din <= x"000a23d9";
		wait for Clk_period;
		Addr <=  "0100011110010";
		Trees_din <= x"ac000704";
		wait for Clk_period;
		Addr <=  "0100011110011";
		Trees_din <= x"007223d9";
		wait for Clk_period;
		Addr <=  "0100011110100";
		Trees_din <= x"002023d9";
		wait for Clk_period;
		Addr <=  "0100011110101";
		Trees_din <= x"ffe723d9";
		wait for Clk_period;
		Addr <=  "0100011110110";
		Trees_din <= x"d2feb620";
		wait for Clk_period;
		Addr <=  "0100011110111";
		Trees_din <= x"dc001e10";
		wait for Clk_period;
		Addr <=  "0100011111000";
		Trees_din <= x"c8ffb208";
		wait for Clk_period;
		Addr <=  "0100011111001";
		Trees_din <= x"10ff6304";
		wait for Clk_period;
		Addr <=  "0100011111010";
		Trees_din <= x"003b248d";
		wait for Clk_period;
		Addr <=  "0100011111011";
		Trees_din <= x"ffc1248d";
		wait for Clk_period;
		Addr <=  "0100011111100";
		Trees_din <= x"d3fe9404";
		wait for Clk_period;
		Addr <=  "0100011111101";
		Trees_din <= x"ffe1248d";
		wait for Clk_period;
		Addr <=  "0100011111110";
		Trees_din <= x"ff86248d";
		wait for Clk_period;
		Addr <=  "0100011111111";
		Trees_din <= x"52ff5b08";
		wait for Clk_period;
		Addr <=  "0100100000000";
		Trees_din <= x"9cffb004";
		wait for Clk_period;
		Addr <=  "0100100000001";
		Trees_din <= x"ffb2248d";
		wait for Clk_period;
		Addr <=  "0100100000010";
		Trees_din <= x"0015248d";
		wait for Clk_period;
		Addr <=  "0100100000011";
		Trees_din <= x"73ffaf04";
		wait for Clk_period;
		Addr <=  "0100100000100";
		Trees_din <= x"0057248d";
		wait for Clk_period;
		Addr <=  "0100100000101";
		Trees_din <= x"0001248d";
		wait for Clk_period;
		Addr <=  "0100100000110";
		Trees_din <= x"53ff751c";
		wait for Clk_period;
		Addr <=  "0100100000111";
		Trees_din <= x"15ff800c";
		wait for Clk_period;
		Addr <=  "0100100001000";
		Trees_din <= x"14ff6d08";
		wait for Clk_period;
		Addr <=  "0100100001001";
		Trees_din <= x"c4fec704";
		wait for Clk_period;
		Addr <=  "0100100001010";
		Trees_din <= x"ffee248d";
		wait for Clk_period;
		Addr <=  "0100100001011";
		Trees_din <= x"ff8d248d";
		wait for Clk_period;
		Addr <=  "0100100001100";
		Trees_din <= x"0006248d";
		wait for Clk_period;
		Addr <=  "0100100001101";
		Trees_din <= x"f1ffae04";
		wait for Clk_period;
		Addr <=  "0100100001110";
		Trees_din <= x"ffbb248d";
		wait for Clk_period;
		Addr <=  "0100100001111";
		Trees_din <= x"c1fedd08";
		wait for Clk_period;
		Addr <=  "0100100010000";
		Trees_din <= x"42ff6204";
		wait for Clk_period;
		Addr <=  "0100100010001";
		Trees_din <= x"fff4248d";
		wait for Clk_period;
		Addr <=  "0100100010010";
		Trees_din <= x"004f248d";
		wait for Clk_period;
		Addr <=  "0100100010011";
		Trees_din <= x"ffdb248d";
		wait for Clk_period;
		Addr <=  "0100100010100";
		Trees_din <= x"f9ff991c";
		wait for Clk_period;
		Addr <=  "0100100010101";
		Trees_din <= x"37ff6010";
		wait for Clk_period;
		Addr <=  "0100100010110";
		Trees_din <= x"3aff2308";
		wait for Clk_period;
		Addr <=  "0100100010111";
		Trees_din <= x"25001304";
		wait for Clk_period;
		Addr <=  "0100100011000";
		Trees_din <= x"0043248d";
		wait for Clk_period;
		Addr <=  "0100100011001";
		Trees_din <= x"ffe6248d";
		wait for Clk_period;
		Addr <=  "0100100011010";
		Trees_din <= x"7bfec704";
		wait for Clk_period;
		Addr <=  "0100100011011";
		Trees_din <= x"000d248d";
		wait for Clk_period;
		Addr <=  "0100100011100";
		Trees_din <= x"ffa8248d";
		wait for Clk_period;
		Addr <=  "0100100011101";
		Trees_din <= x"e5ff3408";
		wait for Clk_period;
		Addr <=  "0100100011110";
		Trees_din <= x"da000104";
		wait for Clk_period;
		Addr <=  "0100100011111";
		Trees_din <= x"005a248d";
		wait for Clk_period;
		Addr <=  "0100100100000";
		Trees_din <= x"fffd248d";
		wait for Clk_period;
		Addr <=  "0100100100001";
		Trees_din <= x"ffd4248d";
		wait for Clk_period;
		Addr <=  "0100100100010";
		Trees_din <= x"ffc1248d";
		wait for Clk_period;
		Addr <=  "0100100100011";
		Trees_din <= x"8dfe4b08";
		wait for Clk_period;
		Addr <=  "0100100100100";
		Trees_din <= x"d1ff6204";
		wait for Clk_period;
		Addr <=  "0100100100101";
		Trees_din <= x"ff9a2531";
		wait for Clk_period;
		Addr <=  "0100100100110";
		Trees_din <= x"00182531";
		wait for Clk_period;
		Addr <=  "0100100100111";
		Trees_din <= x"c4ff0628";
		wait for Clk_period;
		Addr <=  "0100100101000";
		Trees_din <= x"18ffe71c";
		wait for Clk_period;
		Addr <=  "0100100101001";
		Trees_din <= x"24ffe110";
		wait for Clk_period;
		Addr <=  "0100100101010";
		Trees_din <= x"86ff5e08";
		wait for Clk_period;
		Addr <=  "0100100101011";
		Trees_din <= x"34001004";
		wait for Clk_period;
		Addr <=  "0100100101100";
		Trees_din <= x"004e2531";
		wait for Clk_period;
		Addr <=  "0100100101101";
		Trees_din <= x"ffec2531";
		wait for Clk_period;
		Addr <=  "0100100101110";
		Trees_din <= x"41ff2a04";
		wait for Clk_period;
		Addr <=  "0100100101111";
		Trees_din <= x"ffba2531";
		wait for Clk_period;
		Addr <=  "0100100110000";
		Trees_din <= x"000a2531";
		wait for Clk_period;
		Addr <=  "0100100110001";
		Trees_din <= x"3dffc004";
		wait for Clk_period;
		Addr <=  "0100100110010";
		Trees_din <= x"00072531";
		wait for Clk_period;
		Addr <=  "0100100110011";
		Trees_din <= x"7cff6f04";
		wait for Clk_period;
		Addr <=  "0100100110100";
		Trees_din <= x"001f2531";
		wait for Clk_period;
		Addr <=  "0100100110101";
		Trees_din <= x"006d2531";
		wait for Clk_period;
		Addr <=  "0100100110110";
		Trees_din <= x"adff3104";
		wait for Clk_period;
		Addr <=  "0100100110111";
		Trees_din <= x"00342531";
		wait for Clk_period;
		Addr <=  "0100100111000";
		Trees_din <= x"cbff5c04";
		wait for Clk_period;
		Addr <=  "0100100111001";
		Trees_din <= x"00052531";
		wait for Clk_period;
		Addr <=  "0100100111010";
		Trees_din <= x"ff9c2531";
		wait for Clk_period;
		Addr <=  "0100100111011";
		Trees_din <= x"c1fedf18";
		wait for Clk_period;
		Addr <=  "0100100111100";
		Trees_din <= x"d800320c";
		wait for Clk_period;
		Addr <=  "0100100111101";
		Trees_din <= x"57ff7508";
		wait for Clk_period;
		Addr <=  "0100100111110";
		Trees_din <= x"1afea104";
		wait for Clk_period;
		Addr <=  "0100100111111";
		Trees_din <= x"fffa2531";
		wait for Clk_period;
		Addr <=  "0100101000000";
		Trees_din <= x"ff9c2531";
		wait for Clk_period;
		Addr <=  "0100101000001";
		Trees_din <= x"001c2531";
		wait for Clk_period;
		Addr <=  "0100101000010";
		Trees_din <= x"07009a08";
		wait for Clk_period;
		Addr <=  "0100101000011";
		Trees_din <= x"c7ff9f04";
		wait for Clk_period;
		Addr <=  "0100101000100";
		Trees_din <= x"00362531";
		wait for Clk_period;
		Addr <=  "0100101000101";
		Trees_din <= x"ffe12531";
		wait for Clk_period;
		Addr <=  "0100101000110";
		Trees_din <= x"ffbe2531";
		wait for Clk_period;
		Addr <=  "0100101000111";
		Trees_din <= x"b5ff5b04";
		wait for Clk_period;
		Addr <=  "0100101001000";
		Trees_din <= x"ff932531";
		wait for Clk_period;
		Addr <=  "0100101001001";
		Trees_din <= x"06ffe004";
		wait for Clk_period;
		Addr <=  "0100101001010";
		Trees_din <= x"ffdf2531";
		wait for Clk_period;
		Addr <=  "0100101001011";
		Trees_din <= x"003e2531";
		wait for Clk_period;
		Addr <=  "0100101001100";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  3
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"0c001844";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"1400973c";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"32ffa620";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"14ffc510";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"e8007b08";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"c1001f04";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"ff5200bd";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"000f00bd";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"0cffc204";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"ff7400bd";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"01b000bd";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"69feef08";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"53ff7404";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"ff9600bd";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"02e700bd";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"a9fef304";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"002a00bd";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"ff5900bd";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"86fff910";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"13002608";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"f7feef04";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"01cc00bd";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"ffe300bd";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"85001c04";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"ff6200bd";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"003300bd";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"0cff2104";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"ff9c00bd";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"1cffa604";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"038d00bd";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"00ca00bd";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"50ff2f04";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"037a00bd";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"00a600bd";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"ebff6e0c";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"96fff408";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"04ffd704";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"003700bd";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"ff6000bd";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"028200bd";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"8cffc20c";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"83ff9b08";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"96ff3c04";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"015c00bd";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"049b00bd";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"008900bd";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"005b00bd";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"0cffcf44";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"14ffe520";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"95001514";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"9200040c";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"c1001f08";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"0effe904";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"ff580199";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"ffe30199";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"00280199";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"1b003f04";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"ff6f0199";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"01660199";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"b0ffc504";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"ff630199";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"6bff0e04";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"ffa10199";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"02500199";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"53fffe10";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"9dffe10c";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"14006d04";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"ff5d0199";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"87ff7b04";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"ffa40199";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"00d80199";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"00d60199";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"77ff6508";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"5d001e04";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"ff6d0199";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"010c0199";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"64ff4e08";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"19fef504";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"00250199";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"02350199";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"ffa50199";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"ebff6310";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"e8005708";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"2a00db04";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"ff5f0199";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"00390199";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"23ffa204";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"ffa30199";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"01b80199";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"f7ff8910";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"0bffa304";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"fffa0199";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"3aff7008";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"bafff804";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"01d90199";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"00070199";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"00080199";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"94ffbc08";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"16fef704";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"01450199";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"00140199";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"ff780199";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"0cffcf44";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"14ffe524";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"95001518";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"92000410";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"0eff9b08";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"0cffc204";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"ff5b0265";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"fff00265";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"96ff9b04";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"ff640265";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"007c0265";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"baff8904";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"01240265";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"ff740265";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"b0ffc504";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"ff680265";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"6bff3d04";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"ffee0265";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"02090265";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"70ff3d08";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"32ff4604";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"00300265";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"ff610265";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"f3ff3e10";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"8dff2608";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"4dfe5004";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"ffa10265";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"018a0265";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"58fecd04";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"00420265";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"ff870265";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"d000a804";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"ff6e0265";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"00300265";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"ebff6310";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"e8005708";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"3cff8b04";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"ff630265";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"00370265";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"3f004704";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"01430265";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"ffa10265";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"8cffe210";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"15ff4804";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"ff910265";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"97ffb908";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"e9fefd04";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"ffe80265";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"014b0265";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"ff9a0265";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"ff830265";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"0cffcf4c";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"92ffd12c";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"0eff9b1c";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"95001510";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"0cffc208";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"7f009e04";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"ff5e0359";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"fff20359";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"d2ff7504";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"ff900359";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"00cd0359";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"b0ffc504";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"ff6d0359";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"56ff4a04";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"ffa20359";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"01510359";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"4f002d08";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"98ff6304";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"ff660359";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"00c10359";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"2bff1604";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"ffab0359";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"01280359";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"70ff3208";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"3fffd304";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"00860359";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"ff660359";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"f1ffa908";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"78ff2e04";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"00280359";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"ff7b0359";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"96ff7108";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"a7003604";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"ff840359";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"002e0359";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"c1feb504";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"fffd0359";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"01650359";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"ebff6310";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"e8005708";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"a4fed904";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"00380359";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"ff660359";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"45fedf04";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"01060359";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"ffa10359";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"c1fec90c";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"8dfefc08";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"03ffca04";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"00c20359";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"00220359";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"ff610359";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"84ffdc08";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"85000a04";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"ff8a0359";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"00aa0359";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"e9ff0e04";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"ffeb0359";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"bafff804";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"01130359";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"002b0359";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"0cffcf44";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"92ffd128";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"9500151c";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"14ffee10";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"34ffbe08";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"e8006e04";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"ff7b043d";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"0100043d";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"4300c204";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"ff5e043d";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"000e043d";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"77ff8004";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"ff6b043d";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"8dfefe04";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"00ef043d";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"ffab043d";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"6bff1804";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"ff6f043d";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"e0ff7304";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"ff9e043d";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"0135043d";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"70ff3208";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"87feec04";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"0078043d";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"ff6a043d";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"c7ff6208";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"f1000304";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"ff7e043d";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"002d043d";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"64ff6f08";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"ed000704";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"00fb043d";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"ffa4043d";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"ff93043d";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"ebff6310";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"e8005708";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"42001d04";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"ff6a043d";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"0039043d";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"94ff8304";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"ffa3043d";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"00d8043d";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"c1fec90c";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"8dfefc08";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"0fff5404";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"00ae043d";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"0019043d";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"ff67043d";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"15ff4804";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"ffa1043d";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"bafff808";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"84ffdc04";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"0024043d";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"00eb043d";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"16ff8304";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"ff93043d";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"0083043d";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"0cffc250";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"92ffd130";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"0eff9b1c";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"95001510";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"70ff9508";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"7f009e04";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"ff600529";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"001a0529";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"d800a504";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"ff770529";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"00d90529";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"b0ffc504";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"ff770529";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"54004504";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"ffa70529";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"00f60529";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"15ff7d04";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"ff710529";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"96ff8e08";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"31ff0f04";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"00110529";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"ff900529";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"1dff3104";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"013c0529";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"00490529";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"f1ffaa08";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"b7005004";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"ff710529";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"00160529";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"96ff7108";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"7ffef404";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"002b0529";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"ff760529";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"18ff9f08";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"ddff8104";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"ff900529";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"002a0529";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"f2014d04";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"ffce0529";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"01050529";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"ebff6310";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"e8005708";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"5cff2604";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"00370529";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"ff6c0529";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"31ff8b04";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"00b70529";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"ffa20529";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"15ff4804";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"ff890529";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"97ff830c";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"8cffdb08";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"ac008104";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"00d30529";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"000a0529";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"ffe60529";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"0dff3304";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"003e0529";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"ff850529";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"0cffc254";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"92ffd130";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"0eff9b1c";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"95001510";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"70ff9508";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"7f009e04";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"ff620625";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"00170625";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"d800a504";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"ff7c0625";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"00b80625";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"6bff1804";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"ff7a0625";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"b2ffe404";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"ffab0625";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"00db0625";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"15ff7d04";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"ff760625";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"96ff8e08";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"beffa304";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"00120625";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"ff960625";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"1dff3104";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"010e0625";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"003e0625";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"c7ff6208";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"e6ff0404";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"00830625";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"ff700625";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"18ffdf0c";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"dc002a04";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"ff770625";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"06ffe804";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"ffe90625";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"00be0625";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"37ff5b08";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"f1ffa604";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"00100625";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"01160625";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"3bff1004";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"008f0625";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"ff890625";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"e9ff2a0c";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"e7ffc504";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"ff6b0625";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"80ffaf04";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"fff40625";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"007b0625";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"bafff818";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"e8ff9d08";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"d7004204";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"fff10625";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"ff950625";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"c1feb208";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"0fff4404";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"006b0625";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"ff920625";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"72ffa304";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"001c0625";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"00c40625";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"f8ffa404";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"005a0625";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"ff7c0625";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"32ffa640";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"13004620";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"e9ff7b10";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"6f00110c";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"92ffc808";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"b9ffd004";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"ff660719";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"fff60719";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"00430719";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"007f0719";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"12ff9304";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"ff820719";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"9cffba08";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"34ffe904";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"010e0719";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"001d0719";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"ffa40719";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"14ffee18";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"9dfe8408";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"e3fec804";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"ff9c0719";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"00820719";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"1e00c408";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"8100a204";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"ff610719";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"fffb0719";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"16ff1d04";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"ffa50719";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"00420719";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"53ffef04";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"ff8f0719";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"007c0719";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"c0ff7208";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"fbfee104";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"00410719";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"ff6a0719";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"baff8a18";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"31ffad10";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"c2ffb508";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"49ffff04";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"00c70719";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"002d0719";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"27ff6f04";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"004c0719";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"ff9e0719";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"cafed904";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"ff8a0719";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"00450719";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"5fff290c";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"efff2008";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"0bffdc04";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"ffa50719";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"00740719";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"ff580719";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"f1ff8f08";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"d700a804";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"ff8e0719";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"00120719";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"fdffa004";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"00a20719";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"ffca0719";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"32ffa644";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"13004624";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"e9ff7b14";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"e5ff650c";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"a5fe9c08";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"65ff1804";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"00940805";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"ffa70805";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"ff680805";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"98fe4c04";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"00c40805";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"ffa80805";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"12ff9304";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"ff860805";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"cf003f08";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"bcfeff04";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"ffd60805";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"00ec0805";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"ffa70805";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"14ffcf14";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"9dfe8408";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"51ffdf04";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"ffa00805";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"007a0805";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"6f009a04";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"ff620805";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"a0fef304";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"ffae0805";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"00420805";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"63ffd204";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"ff810805";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"71ff6104";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"00920805";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"ffd90805";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"c0ff7208";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"fbfee104";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"00350805";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"ff6d0805";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"c1fec314";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"45febe0c";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"ac003408";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"31ff7204";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"009e0805";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"002c0805";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"ffa60805";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"b6fee304";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"00000805";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"ff690805";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"83ff950c";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"6ffee904";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"ff8b0805";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"15ff5304";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"000a0805";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"00af0805";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"8affb704";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"ff720805";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"60ffb704";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"000a0805";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"007f0805";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"32ffa644";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"13004628";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"ebff4414";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"e3ff5510";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"95ffff08";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"2e005904";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"ff6a0901";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"ffe90901";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"feffa004";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"ffad0901";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"00880901";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"00910901";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"52ff180c";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"cf003f08";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"d8005f04";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"00130901";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"00f60901";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"ffd50901";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"81000004";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"ff8e0901";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"00160901";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"14ffcf10";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"4cfe1004";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"00250901";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"1e00c408";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"4f013d04";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"ff630901";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"ffce0901";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"fffc0901";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"e4ff1b04";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"ff840901";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"00ff9304";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"ffd80901";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"008d0901";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"c0ff7208";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"52feca04";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"00340901";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"ff700901";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"baff8a18";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"31ffad10";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"49ffff08";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"c2ffb504";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"00b30901";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"fff80901";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"f1000f04";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"ffa80901";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"00720901";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"cafed904";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"ff930901";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"00360901";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"73ffd90c";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"0bffc604";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"ff950901";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"27ff8c04";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"000f0901";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"00ae0901";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"faffcb08";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"a7fff704";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"ff630901";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"00390901";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"f0ff6904";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"00780901";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"00090901";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"32ffa648";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"1300462c";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"3cfec210";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"e8000c04";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"ff9e0a01";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"9affd604";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"fff10a01";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"27ff9004";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"013b0a01";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"004e0a01";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"ebff560c";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"0cffcf04";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"ff6c0a01";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"1effcb04";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"ffd20a01";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"00570a01";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"c2ff1e08";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"d9ffde04";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"000c0a01";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"009d0a01";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"b6ff3b04";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"000d0a01";
		wait for Clk_period;
		Addr <=  "0001001010111";
		Trees_din <= x"ff9b0a01";
		wait for Clk_period;
		Addr <=  "0001001011000";
		Trees_din <= x"b1fffb14";
		wait for Clk_period;
		Addr <=  "0001001011001";
		Trees_din <= x"14ffcf0c";
		wait for Clk_period;
		Addr <=  "0001001011010";
		Trees_din <= x"6f009a08";
		wait for Clk_period;
		Addr <=  "0001001011011";
		Trees_din <= x"4f013d04";
		wait for Clk_period;
		Addr <=  "0001001011100";
		Trees_din <= x"ff640a01";
		wait for Clk_period;
		Addr <=  "0001001011101";
		Trees_din <= x"ffd70a01";
		wait for Clk_period;
		Addr <=  "0001001011110";
		Trees_din <= x"000a0a01";
		wait for Clk_period;
		Addr <=  "0001001011111";
		Trees_din <= x"2fffcf04";
		wait for Clk_period;
		Addr <=  "0001001100000";
		Trees_din <= x"ff930a01";
		wait for Clk_period;
		Addr <=  "0001001100001";
		Trees_din <= x"00660a01";
		wait for Clk_period;
		Addr <=  "0001001100010";
		Trees_din <= x"e4ff0904";
		wait for Clk_period;
		Addr <=  "0001001100011";
		Trees_din <= x"ff9e0a01";
		wait for Clk_period;
		Addr <=  "0001001100100";
		Trees_din <= x"00ae0a01";
		wait for Clk_period;
		Addr <=  "0001001100101";
		Trees_din <= x"c0ff7208";
		wait for Clk_period;
		Addr <=  "0001001100110";
		Trees_din <= x"52feca04";
		wait for Clk_period;
		Addr <=  "0001001100111";
		Trees_din <= x"002e0a01";
		wait for Clk_period;
		Addr <=  "0001001101000";
		Trees_din <= x"ff740a01";
		wait for Clk_period;
		Addr <=  "0001001101001";
		Trees_din <= x"baff6714";
		wait for Clk_period;
		Addr <=  "0001001101010";
		Trees_din <= x"cbff8404";
		wait for Clk_period;
		Addr <=  "0001001101011";
		Trees_din <= x"ff9b0a01";
		wait for Clk_period;
		Addr <=  "0001001101100";
		Trees_din <= x"70ff1008";
		wait for Clk_period;
		Addr <=  "0001001101101";
		Trees_din <= x"0a011804";
		wait for Clk_period;
		Addr <=  "0001001101110";
		Trees_din <= x"ff920a01";
		wait for Clk_period;
		Addr <=  "0001001101111";
		Trees_din <= x"00710a01";
		wait for Clk_period;
		Addr <=  "0001001110000";
		Trees_din <= x"15ff2d04";
		wait for Clk_period;
		Addr <=  "0001001110001";
		Trees_din <= x"00100a01";
		wait for Clk_period;
		Addr <=  "0001001110010";
		Trees_din <= x"00b40a01";
		wait for Clk_period;
		Addr <=  "0001001110011";
		Trees_din <= x"f1ff9e0c";
		wait for Clk_period;
		Addr <=  "0001001110100";
		Trees_din <= x"fbff3708";
		wait for Clk_period;
		Addr <=  "0001001110101";
		Trees_din <= x"3bff2604";
		wait for Clk_period;
		Addr <=  "0001001110110";
		Trees_din <= x"00660a01";
		wait for Clk_period;
		Addr <=  "0001001110111";
		Trees_din <= x"ffe70a01";
		wait for Clk_period;
		Addr <=  "0001001111000";
		Trees_din <= x"ff760a01";
		wait for Clk_period;
		Addr <=  "0001001111001";
		Trees_din <= x"27ff5f08";
		wait for Clk_period;
		Addr <=  "0001001111010";
		Trees_din <= x"51fffc04";
		wait for Clk_period;
		Addr <=  "0001001111011";
		Trees_din <= x"ff710a01";
		wait for Clk_period;
		Addr <=  "0001001111100";
		Trees_din <= x"005a0a01";
		wait for Clk_period;
		Addr <=  "0001001111101";
		Trees_din <= x"96ff6504";
		wait for Clk_period;
		Addr <=  "0001001111110";
		Trees_din <= x"ffba0a01";
		wait for Clk_period;
		Addr <=  "0001001111111";
		Trees_din <= x"00970a01";
		wait for Clk_period;
		Addr <=  "0001010000000";
		Trees_din <= x"32ff973c";
		wait for Clk_period;
		Addr <=  "0001010000001";
		Trees_din <= x"13004624";
		wait for Clk_period;
		Addr <=  "0001010000010";
		Trees_din <= x"d4ff770c";
		wait for Clk_period;
		Addr <=  "0001010000011";
		Trees_din <= x"f4ffb304";
		wait for Clk_period;
		Addr <=  "0001010000100";
		Trees_din <= x"ff6f0aed";
		wait for Clk_period;
		Addr <=  "0001010000101";
		Trees_din <= x"6affa004";
		wait for Clk_period;
		Addr <=  "0001010000110";
		Trees_din <= x"ffe20aed";
		wait for Clk_period;
		Addr <=  "0001010000111";
		Trees_din <= x"005f0aed";
		wait for Clk_period;
		Addr <=  "0001010001000";
		Trees_din <= x"e8000508";
		wait for Clk_period;
		Addr <=  "0001010001001";
		Trees_din <= x"9ffef304";
		wait for Clk_period;
		Addr <=  "0001010001010";
		Trees_din <= x"001e0aed";
		wait for Clk_period;
		Addr <=  "0001010001011";
		Trees_din <= x"ff8a0aed";
		wait for Clk_period;
		Addr <=  "0001010001100";
		Trees_din <= x"3cfec208";
		wait for Clk_period;
		Addr <=  "0001010001101";
		Trees_din <= x"14ff4e04";
		wait for Clk_period;
		Addr <=  "0001010001110";
		Trees_din <= x"001f0aed";
		wait for Clk_period;
		Addr <=  "0001010001111";
		Trees_din <= x"01050aed";
		wait for Clk_period;
		Addr <=  "0001010010000";
		Trees_din <= x"86ffba04";
		wait for Clk_period;
		Addr <=  "0001010010001";
		Trees_din <= x"ffae0aed";
		wait for Clk_period;
		Addr <=  "0001010010010";
		Trees_din <= x"00720aed";
		wait for Clk_period;
		Addr <=  "0001010010011";
		Trees_din <= x"b1fffb10";
		wait for Clk_period;
		Addr <=  "0001010010100";
		Trees_din <= x"1e00c40c";
		wait for Clk_period;
		Addr <=  "0001010010101";
		Trees_din <= x"a3fe6e04";
		wait for Clk_period;
		Addr <=  "0001010010110";
		Trees_din <= x"fffa0aed";
		wait for Clk_period;
		Addr <=  "0001010010111";
		Trees_din <= x"2b014504";
		wait for Clk_period;
		Addr <=  "0001010011000";
		Trees_din <= x"ff650aed";
		wait for Clk_period;
		Addr <=  "0001010011001";
		Trees_din <= x"ffce0aed";
		wait for Clk_period;
		Addr <=  "0001010011010";
		Trees_din <= x"00130aed";
		wait for Clk_period;
		Addr <=  "0001010011011";
		Trees_din <= x"e4ff0904";
		wait for Clk_period;
		Addr <=  "0001010011100";
		Trees_din <= x"ffa40aed";
		wait for Clk_period;
		Addr <=  "0001010011101";
		Trees_din <= x"009e0aed";
		wait for Clk_period;
		Addr <=  "0001010011110";
		Trees_din <= x"0cff1c10";
		wait for Clk_period;
		Addr <=  "0001010011111";
		Trees_din <= x"13001b08";
		wait for Clk_period;
		Addr <=  "0001010100000";
		Trees_din <= x"efff7b04";
		wait for Clk_period;
		Addr <=  "0001010100001";
		Trees_din <= x"ff9e0aed";
		wait for Clk_period;
		Addr <=  "0001010100010";
		Trees_din <= x"00b50aed";
		wait for Clk_period;
		Addr <=  "0001010100011";
		Trees_din <= x"9cfecf04";
		wait for Clk_period;
		Addr <=  "0001010100100";
		Trees_din <= x"ffec0aed";
		wait for Clk_period;
		Addr <=  "0001010100101";
		Trees_din <= x"ff710aed";
		wait for Clk_period;
		Addr <=  "0001010100110";
		Trees_din <= x"baff7410";
		wait for Clk_period;
		Addr <=  "0001010100111";
		Trees_din <= x"1effe90c";
		wait for Clk_period;
		Addr <=  "0001010101000";
		Trees_din <= x"97ff9308";
		wait for Clk_period;
		Addr <=  "0001010101001";
		Trees_din <= x"31ffad04";
		wait for Clk_period;
		Addr <=  "0001010101010";
		Trees_din <= x"00a90aed";
		wait for Clk_period;
		Addr <=  "0001010101011";
		Trees_din <= x"ffff0aed";
		wait for Clk_period;
		Addr <=  "0001010101100";
		Trees_din <= x"ffd00aed";
		wait for Clk_period;
		Addr <=  "0001010101101";
		Trees_din <= x"ffd90aed";
		wait for Clk_period;
		Addr <=  "0001010101110";
		Trees_din <= x"dfff1c0c";
		wait for Clk_period;
		Addr <=  "0001010101111";
		Trees_din <= x"b3ff6f08";
		wait for Clk_period;
		Addr <=  "0001010110000";
		Trees_din <= x"96ff9f04";
		wait for Clk_period;
		Addr <=  "0001010110001";
		Trees_din <= x"001f0aed";
		wait for Clk_period;
		Addr <=  "0001010110010";
		Trees_din <= x"009e0aed";
		wait for Clk_period;
		Addr <=  "0001010110011";
		Trees_din <= x"ffcb0aed";
		wait for Clk_period;
		Addr <=  "0001010110100";
		Trees_din <= x"51000208";
		wait for Clk_period;
		Addr <=  "0001010110101";
		Trees_din <= x"97feb704";
		wait for Clk_period;
		Addr <=  "0001010110110";
		Trees_din <= x"00450aed";
		wait for Clk_period;
		Addr <=  "0001010110111";
		Trees_din <= x"ff810aed";
		wait for Clk_period;
		Addr <=  "0001010111000";
		Trees_din <= x"a3ff1d04";
		wait for Clk_period;
		Addr <=  "0001010111001";
		Trees_din <= x"008f0aed";
		wait for Clk_period;
		Addr <=  "0001010111010";
		Trees_din <= x"ffbe0aed";
		wait for Clk_period;
		Addr <=  "0001010111011";
		Trees_din <= x"32ff9738";
		wait for Clk_period;
		Addr <=  "0001010111100";
		Trees_din <= x"13004620";
		wait for Clk_period;
		Addr <=  "0001010111101";
		Trees_din <= x"d4ff7708";
		wait for Clk_period;
		Addr <=  "0001010111110";
		Trees_din <= x"f4ffb304";
		wait for Clk_period;
		Addr <=  "0001010111111";
		Trees_din <= x"ff710bc1";
		wait for Clk_period;
		Addr <=  "0001011000000";
		Trees_din <= x"002a0bc1";
		wait for Clk_period;
		Addr <=  "0001011000001";
		Trees_din <= x"e8000508";
		wait for Clk_period;
		Addr <=  "0001011000010";
		Trees_din <= x"4dfef904";
		wait for Clk_period;
		Addr <=  "0001011000011";
		Trees_din <= x"ff8e0bc1";
		wait for Clk_period;
		Addr <=  "0001011000100";
		Trees_din <= x"001f0bc1";
		wait for Clk_period;
		Addr <=  "0001011000101";
		Trees_din <= x"d2ff0b08";
		wait for Clk_period;
		Addr <=  "0001011000110";
		Trees_din <= x"0eff4704";
		wait for Clk_period;
		Addr <=  "0001011000111";
		Trees_din <= x"ffa90bc1";
		wait for Clk_period;
		Addr <=  "0001011001000";
		Trees_din <= x"00340bc1";
		wait for Clk_period;
		Addr <=  "0001011001001";
		Trees_din <= x"34ffe904";
		wait for Clk_period;
		Addr <=  "0001011001010";
		Trees_din <= x"00d20bc1";
		wait for Clk_period;
		Addr <=  "0001011001011";
		Trees_din <= x"001c0bc1";
		wait for Clk_period;
		Addr <=  "0001011001100";
		Trees_din <= x"b1fffb10";
		wait for Clk_period;
		Addr <=  "0001011001101";
		Trees_din <= x"6f009a0c";
		wait for Clk_period;
		Addr <=  "0001011001110";
		Trees_din <= x"a3fe6e04";
		wait for Clk_period;
		Addr <=  "0001011001111";
		Trees_din <= x"fffb0bc1";
		wait for Clk_period;
		Addr <=  "0001011010000";
		Trees_din <= x"2b014504";
		wait for Clk_period;
		Addr <=  "0001011010001";
		Trees_din <= x"ff650bc1";
		wait for Clk_period;
		Addr <=  "0001011010010";
		Trees_din <= x"ffd00bc1";
		wait for Clk_period;
		Addr <=  "0001011010011";
		Trees_din <= x"001d0bc1";
		wait for Clk_period;
		Addr <=  "0001011010100";
		Trees_din <= x"63ffe904";
		wait for Clk_period;
		Addr <=  "0001011010101";
		Trees_din <= x"ffa80bc1";
		wait for Clk_period;
		Addr <=  "0001011010110";
		Trees_din <= x"00930bc1";
		wait for Clk_period;
		Addr <=  "0001011010111";
		Trees_din <= x"c0ff6408";
		wait for Clk_period;
		Addr <=  "0001011011000";
		Trees_din <= x"fdff0304";
		wait for Clk_period;
		Addr <=  "0001011011001";
		Trees_din <= x"ffe60bc1";
		wait for Clk_period;
		Addr <=  "0001011011010";
		Trees_din <= x"ff7a0bc1";
		wait for Clk_period;
		Addr <=  "0001011011011";
		Trees_din <= x"c1feb30c";
		wait for Clk_period;
		Addr <=  "0001011011100";
		Trees_din <= x"18003d08";
		wait for Clk_period;
		Addr <=  "0001011011101";
		Trees_din <= x"01fe6304";
		wait for Clk_period;
		Addr <=  "0001011011110";
		Trees_din <= x"ffe90bc1";
		wait for Clk_period;
		Addr <=  "0001011011111";
		Trees_din <= x"ff7f0bc1";
		wait for Clk_period;
		Addr <=  "0001011100000";
		Trees_din <= x"00270bc1";
		wait for Clk_period;
		Addr <=  "0001011100001";
		Trees_din <= x"83ff7110";
		wait for Clk_period;
		Addr <=  "0001011100010";
		Trees_din <= x"f1ff9008";
		wait for Clk_period;
		Addr <=  "0001011100011";
		Trees_din <= x"baff6704";
		wait for Clk_period;
		Addr <=  "0001011100100";
		Trees_din <= x"006f0bc1";
		wait for Clk_period;
		Addr <=  "0001011100101";
		Trees_din <= x"ffb30bc1";
		wait for Clk_period;
		Addr <=  "0001011100110";
		Trees_din <= x"a6ffa704";
		wait for Clk_period;
		Addr <=  "0001011100111";
		Trees_din <= x"009a0bc1";
		wait for Clk_period;
		Addr <=  "0001011101000";
		Trees_din <= x"ffce0bc1";
		wait for Clk_period;
		Addr <=  "0001011101001";
		Trees_din <= x"8affb708";
		wait for Clk_period;
		Addr <=  "0001011101010";
		Trees_din <= x"16ff6e04";
		wait for Clk_period;
		Addr <=  "0001011101011";
		Trees_din <= x"ff730bc1";
		wait for Clk_period;
		Addr <=  "0001011101100";
		Trees_din <= x"ffec0bc1";
		wait for Clk_period;
		Addr <=  "0001011101101";
		Trees_din <= x"8dfee404";
		wait for Clk_period;
		Addr <=  "0001011101110";
		Trees_din <= x"00750bc1";
		wait for Clk_period;
		Addr <=  "0001011101111";
		Trees_din <= x"ffd90bc1";
		wait for Clk_period;
		Addr <=  "0001011110000";
		Trees_din <= x"32ff6e28";
		wait for Clk_period;
		Addr <=  "0001011110001";
		Trees_din <= x"0eff7018";
		wait for Clk_period;
		Addr <=  "0001011110010";
		Trees_din <= x"e8005b0c";
		wait for Clk_period;
		Addr <=  "0001011110011";
		Trees_din <= x"e9001208";
		wait for Clk_period;
		Addr <=  "0001011110100";
		Trees_din <= x"ebffb004";
		wait for Clk_period;
		Addr <=  "0001011110101";
		Trees_din <= x"ff660c85";
		wait for Clk_period;
		Addr <=  "0001011110110";
		Trees_din <= x"ffe90c85";
		wait for Clk_period;
		Addr <=  "0001011110111";
		Trees_din <= x"fff90c85";
		wait for Clk_period;
		Addr <=  "0001011111000";
		Trees_din <= x"d8008f04";
		wait for Clk_period;
		Addr <=  "0001011111001";
		Trees_din <= x"ff870c85";
		wait for Clk_period;
		Addr <=  "0001011111010";
		Trees_din <= x"71ffbd04";
		wait for Clk_period;
		Addr <=  "0001011111011";
		Trees_din <= x"00190c85";
		wait for Clk_period;
		Addr <=  "0001011111100";
		Trees_din <= x"008d0c85";
		wait for Clk_period;
		Addr <=  "0001011111101";
		Trees_din <= x"34ffd608";
		wait for Clk_period;
		Addr <=  "0001011111110";
		Trees_din <= x"3f000004";
		wait for Clk_period;
		Addr <=  "0001011111111";
		Trees_din <= x"00fd0c85";
		wait for Clk_period;
		Addr <=  "0001100000000";
		Trees_din <= x"fffd0c85";
		wait for Clk_period;
		Addr <=  "0001100000001";
		Trees_din <= x"4aff8604";
		wait for Clk_period;
		Addr <=  "0001100000010";
		Trees_din <= x"ff840c85";
		wait for Clk_period;
		Addr <=  "0001100000011";
		Trees_din <= x"00070c85";
		wait for Clk_period;
		Addr <=  "0001100000100";
		Trees_din <= x"0cff1c14";
		wait for Clk_period;
		Addr <=  "0001100000101";
		Trees_din <= x"0dffcd08";
		wait for Clk_period;
		Addr <=  "0001100000110";
		Trees_din <= x"1efee604";
		wait for Clk_period;
		Addr <=  "0001100000111";
		Trees_din <= x"00090c85";
		wait for Clk_period;
		Addr <=  "0001100001000";
		Trees_din <= x"ff730c85";
		wait for Clk_period;
		Addr <=  "0001100001001";
		Trees_din <= x"13004008";
		wait for Clk_period;
		Addr <=  "0001100001010";
		Trees_din <= x"6aff5e04";
		wait for Clk_period;
		Addr <=  "0001100001011";
		Trees_din <= x"00c80c85";
		wait for Clk_period;
		Addr <=  "0001100001100";
		Trees_din <= x"00270c85";
		wait for Clk_period;
		Addr <=  "0001100001101";
		Trees_din <= x"ff9b0c85";
		wait for Clk_period;
		Addr <=  "0001100001110";
		Trees_din <= x"c1feb308";
		wait for Clk_period;
		Addr <=  "0001100001111";
		Trees_din <= x"da005304";
		wait for Clk_period;
		Addr <=  "0001100010000";
		Trees_din <= x"ff810c85";
		wait for Clk_period;
		Addr <=  "0001100010001";
		Trees_din <= x"00240c85";
		wait for Clk_period;
		Addr <=  "0001100010010";
		Trees_din <= x"83ff7110";
		wait for Clk_period;
		Addr <=  "0001100010011";
		Trees_din <= x"baff7608";
		wait for Clk_period;
		Addr <=  "0001100010100";
		Trees_din <= x"f3fe4004";
		wait for Clk_period;
		Addr <=  "0001100010101";
		Trees_din <= x"00000c85";
		wait for Clk_period;
		Addr <=  "0001100010110";
		Trees_din <= x"00a50c85";
		wait for Clk_period;
		Addr <=  "0001100010111";
		Trees_din <= x"0c001804";
		wait for Clk_period;
		Addr <=  "0001100011000";
		Trees_din <= x"ffdd0c85";
		wait for Clk_period;
		Addr <=  "0001100011001";
		Trees_din <= x"00790c85";
		wait for Clk_period;
		Addr <=  "0001100011010";
		Trees_din <= x"8dfee408";
		wait for Clk_period;
		Addr <=  "0001100011011";
		Trees_din <= x"5effeb04";
		wait for Clk_period;
		Addr <=  "0001100011100";
		Trees_din <= x"ffde0c85";
		wait for Clk_period;
		Addr <=  "0001100011101";
		Trees_din <= x"00700c85";
		wait for Clk_period;
		Addr <=  "0001100011110";
		Trees_din <= x"97ff2f04";
		wait for Clk_period;
		Addr <=  "0001100011111";
		Trees_din <= x"ff7d0c85";
		wait for Clk_period;
		Addr <=  "0001100100000";
		Trees_din <= x"00040c85";
		wait for Clk_period;
		Addr <=  "0001100100001";
		Trees_din <= x"14ff4a18";
		wait for Clk_period;
		Addr <=  "0001100100010";
		Trees_din <= x"9dfeb308";
		wait for Clk_period;
		Addr <=  "0001100100011";
		Trees_din <= x"34ffc804";
		wait for Clk_period;
		Addr <=  "0001100100100";
		Trees_din <= x"00a40d49";
		wait for Clk_period;
		Addr <=  "0001100100101";
		Trees_din <= x"ffa30d49";
		wait for Clk_period;
		Addr <=  "0001100100110";
		Trees_din <= x"e3ff6808";
		wait for Clk_period;
		Addr <=  "0001100100111";
		Trees_din <= x"80005904";
		wait for Clk_period;
		Addr <=  "0001100101000";
		Trees_din <= x"ff680d49";
		wait for Clk_period;
		Addr <=  "0001100101001";
		Trees_din <= x"ffd70d49";
		wait for Clk_period;
		Addr <=  "0001100101010";
		Trees_din <= x"0fff3604";
		wait for Clk_period;
		Addr <=  "0001100101011";
		Trees_din <= x"001e0d49";
		wait for Clk_period;
		Addr <=  "0001100101100";
		Trees_din <= x"ffc70d49";
		wait for Clk_period;
		Addr <=  "0001100101101";
		Trees_din <= x"13004f30";
		wait for Clk_period;
		Addr <=  "0001100101110";
		Trees_din <= x"96ffb418";
		wait for Clk_period;
		Addr <=  "0001100101111";
		Trees_din <= x"15ff7608";
		wait for Clk_period;
		Addr <=  "0001100110000";
		Trees_din <= x"7aff1f04";
		wait for Clk_period;
		Addr <=  "0001100110001";
		Trees_din <= x"fff00d49";
		wait for Clk_period;
		Addr <=  "0001100110010";
		Trees_din <= x"ff840d49";
		wait for Clk_period;
		Addr <=  "0001100110011";
		Trees_din <= x"afff8b08";
		wait for Clk_period;
		Addr <=  "0001100110100";
		Trees_din <= x"8cff2304";
		wait for Clk_period;
		Addr <=  "0001100110101";
		Trees_din <= x"003c0d49";
		wait for Clk_period;
		Addr <=  "0001100110110";
		Trees_din <= x"ff8f0d49";
		wait for Clk_period;
		Addr <=  "0001100110111";
		Trees_din <= x"ebff3c04";
		wait for Clk_period;
		Addr <=  "0001100111000";
		Trees_din <= x"ffb00d49";
		wait for Clk_period;
		Addr <=  "0001100111001";
		Trees_din <= x"00980d49";
		wait for Clk_period;
		Addr <=  "0001100111010";
		Trees_din <= x"f9ff6510";
		wait for Clk_period;
		Addr <=  "0001100111011";
		Trees_din <= x"77ff5108";
		wait for Clk_period;
		Addr <=  "0001100111100";
		Trees_din <= x"c1fed904";
		wait for Clk_period;
		Addr <=  "0001100111101";
		Trees_din <= x"ff960d49";
		wait for Clk_period;
		Addr <=  "0001100111110";
		Trees_din <= x"006b0d49";
		wait for Clk_period;
		Addr <=  "0001100111111";
		Trees_din <= x"5bff8c04";
		wait for Clk_period;
		Addr <=  "0001101000000";
		Trees_din <= x"00af0d49";
		wait for Clk_period;
		Addr <=  "0001101000001";
		Trees_din <= x"001c0d49";
		wait for Clk_period;
		Addr <=  "0001101000010";
		Trees_din <= x"f1ffa504";
		wait for Clk_period;
		Addr <=  "0001101000011";
		Trees_din <= x"ffa20d49";
		wait for Clk_period;
		Addr <=  "0001101000100";
		Trees_din <= x"000f0d49";
		wait for Clk_period;
		Addr <=  "0001101000101";
		Trees_din <= x"0cff3d0c";
		wait for Clk_period;
		Addr <=  "0001101000110";
		Trees_din <= x"0eff9b08";
		wait for Clk_period;
		Addr <=  "0001101000111";
		Trees_din <= x"51007304";
		wait for Clk_period;
		Addr <=  "0001101001000";
		Trees_din <= x"ff6d0d49";
		wait for Clk_period;
		Addr <=  "0001101001001";
		Trees_din <= x"ffdc0d49";
		wait for Clk_period;
		Addr <=  "0001101001010";
		Trees_din <= x"002c0d49";
		wait for Clk_period;
		Addr <=  "0001101001011";
		Trees_din <= x"63ff9f04";
		wait for Clk_period;
		Addr <=  "0001101001100";
		Trees_din <= x"ff940d49";
		wait for Clk_period;
		Addr <=  "0001101001101";
		Trees_din <= x"bbff9b08";
		wait for Clk_period;
		Addr <=  "0001101001110";
		Trees_din <= x"c1feb604";
		wait for Clk_period;
		Addr <=  "0001101001111";
		Trees_din <= x"ffcb0d49";
		wait for Clk_period;
		Addr <=  "0001101010000";
		Trees_din <= x"00780d49";
		wait for Clk_period;
		Addr <=  "0001101010001";
		Trees_din <= x"ffa10d49";
		wait for Clk_period;
		Addr <=  "0001101010010";
		Trees_din <= x"14ff4a14";
		wait for Clk_period;
		Addr <=  "0001101010011";
		Trees_din <= x"9dfeb308";
		wait for Clk_period;
		Addr <=  "0001101010100";
		Trees_din <= x"34ffc804";
		wait for Clk_period;
		Addr <=  "0001101010101";
		Trees_din <= x"00930e0d";
		wait for Clk_period;
		Addr <=  "0001101010110";
		Trees_din <= x"ffa80e0d";
		wait for Clk_period;
		Addr <=  "0001101010111";
		Trees_din <= x"e3ff6808";
		wait for Clk_period;
		Addr <=  "0001101011000";
		Trees_din <= x"e9ffe204";
		wait for Clk_period;
		Addr <=  "0001101011001";
		Trees_din <= x"ff680e0d";
		wait for Clk_period;
		Addr <=  "0001101011010";
		Trees_din <= x"ffca0e0d";
		wait for Clk_period;
		Addr <=  "0001101011011";
		Trees_din <= x"fff00e0d";
		wait for Clk_period;
		Addr <=  "0001101011100";
		Trees_din <= x"13004f34";
		wait for Clk_period;
		Addr <=  "0001101011101";
		Trees_din <= x"85fff318";
		wait for Clk_period;
		Addr <=  "0001101011110";
		Trees_din <= x"18001f10";
		wait for Clk_period;
		Addr <=  "0001101011111";
		Trees_din <= x"89fff008";
		wait for Clk_period;
		Addr <=  "0001101100000";
		Trees_din <= x"0c007b04";
		wait for Clk_period;
		Addr <=  "0001101100001";
		Trees_din <= x"ff800e0d";
		wait for Clk_period;
		Addr <=  "0001101100010";
		Trees_din <= x"00110e0d";
		wait for Clk_period;
		Addr <=  "0001101100011";
		Trees_din <= x"4cff5704";
		wait for Clk_period;
		Addr <=  "0001101100100";
		Trees_din <= x"ffc80e0d";
		wait for Clk_period;
		Addr <=  "0001101100101";
		Trees_din <= x"00660e0d";
		wait for Clk_period;
		Addr <=  "0001101100110";
		Trees_din <= x"99feca04";
		wait for Clk_period;
		Addr <=  "0001101100111";
		Trees_din <= x"00950e0d";
		wait for Clk_period;
		Addr <=  "0001101101000";
		Trees_din <= x"ffef0e0d";
		wait for Clk_period;
		Addr <=  "0001101101001";
		Trees_din <= x"03ff630c";
		wait for Clk_period;
		Addr <=  "0001101101010";
		Trees_din <= x"96ff6b08";
		wait for Clk_period;
		Addr <=  "0001101101011";
		Trees_din <= x"29002e04";
		wait for Clk_period;
		Addr <=  "0001101101100";
		Trees_din <= x"ffd10e0d";
		wait for Clk_period;
		Addr <=  "0001101101101";
		Trees_din <= x"006c0e0d";
		wait for Clk_period;
		Addr <=  "0001101101110";
		Trees_din <= x"00a60e0d";
		wait for Clk_period;
		Addr <=  "0001101101111";
		Trees_din <= x"29001c08";
		wait for Clk_period;
		Addr <=  "0001101110000";
		Trees_din <= x"52feef04";
		wait for Clk_period;
		Addr <=  "0001101110001";
		Trees_din <= x"00320e0d";
		wait for Clk_period;
		Addr <=  "0001101110010";
		Trees_din <= x"ff900e0d";
		wait for Clk_period;
		Addr <=  "0001101110011";
		Trees_din <= x"0b00a104";
		wait for Clk_period;
		Addr <=  "0001101110100";
		Trees_din <= x"007e0e0d";
		wait for Clk_period;
		Addr <=  "0001101110101";
		Trees_din <= x"00000e0d";
		wait for Clk_period;
		Addr <=  "0001101110110";
		Trees_din <= x"0cfed404";
		wait for Clk_period;
		Addr <=  "0001101110111";
		Trees_din <= x"ff720e0d";
		wait for Clk_period;
		Addr <=  "0001101111000";
		Trees_din <= x"0eff0e08";
		wait for Clk_period;
		Addr <=  "0001101111001";
		Trees_din <= x"b7002f04";
		wait for Clk_period;
		Addr <=  "0001101111010";
		Trees_din <= x"ff7e0e0d";
		wait for Clk_period;
		Addr <=  "0001101111011";
		Trees_din <= x"000c0e0d";
		wait for Clk_period;
		Addr <=  "0001101111100";
		Trees_din <= x"57ff4e08";
		wait for Clk_period;
		Addr <=  "0001101111101";
		Trees_din <= x"baffa504";
		wait for Clk_period;
		Addr <=  "0001101111110";
		Trees_din <= x"007c0e0d";
		wait for Clk_period;
		Addr <=  "0001101111111";
		Trees_din <= x"ffdc0e0d";
		wait for Clk_period;
		Addr <=  "0001110000000";
		Trees_din <= x"fbfed604";
		wait for Clk_period;
		Addr <=  "0001110000001";
		Trees_din <= x"00020e0d";
		wait for Clk_period;
		Addr <=  "0001110000010";
		Trees_din <= x"ff8f0e0d";
		wait for Clk_period;
		Addr <=  "0001110000011";
		Trees_din <= x"14ff4a14";
		wait for Clk_period;
		Addr <=  "0001110000100";
		Trees_din <= x"9dfeb308";
		wait for Clk_period;
		Addr <=  "0001110000101";
		Trees_din <= x"34ffc804";
		wait for Clk_period;
		Addr <=  "0001110000110";
		Trees_din <= x"008a0ec9";
		wait for Clk_period;
		Addr <=  "0001110000111";
		Trees_din <= x"ffad0ec9";
		wait for Clk_period;
		Addr <=  "0001110001000";
		Trees_din <= x"e3ff6808";
		wait for Clk_period;
		Addr <=  "0001110001001";
		Trees_din <= x"e9ffe204";
		wait for Clk_period;
		Addr <=  "0001110001010";
		Trees_din <= x"ff680ec9";
		wait for Clk_period;
		Addr <=  "0001110001011";
		Trees_din <= x"ffcf0ec9";
		wait for Clk_period;
		Addr <=  "0001110001100";
		Trees_din <= x"fff10ec9";
		wait for Clk_period;
		Addr <=  "0001110001101";
		Trees_din <= x"13004f2c";
		wait for Clk_period;
		Addr <=  "0001110001110";
		Trees_din <= x"96ffb418";
		wait for Clk_period;
		Addr <=  "0001110001111";
		Trees_din <= x"15ff7608";
		wait for Clk_period;
		Addr <=  "0001110010000";
		Trees_din <= x"15ff0904";
		wait for Clk_period;
		Addr <=  "0001110010001";
		Trees_din <= x"ffeb0ec9";
		wait for Clk_period;
		Addr <=  "0001110010010";
		Trees_din <= x"ff8c0ec9";
		wait for Clk_period;
		Addr <=  "0001110010011";
		Trees_din <= x"afffb208";
		wait for Clk_period;
		Addr <=  "0001110010100";
		Trees_din <= x"0cffcf04";
		wait for Clk_period;
		Addr <=  "0001110010101";
		Trees_din <= x"ff9d0ec9";
		wait for Clk_period;
		Addr <=  "0001110010110";
		Trees_din <= x"00210ec9";
		wait for Clk_period;
		Addr <=  "0001110010111";
		Trees_din <= x"70ff5404";
		wait for Clk_period;
		Addr <=  "0001110011000";
		Trees_din <= x"00050ec9";
		wait for Clk_period;
		Addr <=  "0001110011001";
		Trees_din <= x"008b0ec9";
		wait for Clk_period;
		Addr <=  "0001110011010";
		Trees_din <= x"f9ff6510";
		wait for Clk_period;
		Addr <=  "0001110011011";
		Trees_din <= x"e5fe8c08";
		wait for Clk_period;
		Addr <=  "0001110011100";
		Trees_din <= x"f7ff4404";
		wait for Clk_period;
		Addr <=  "0001110011101";
		Trees_din <= x"00520ec9";
		wait for Clk_period;
		Addr <=  "0001110011110";
		Trees_din <= x"ffb20ec9";
		wait for Clk_period;
		Addr <=  "0001110011111";
		Trees_din <= x"5bff8c04";
		wait for Clk_period;
		Addr <=  "0001110100000";
		Trees_din <= x"009e0ec9";
		wait for Clk_period;
		Addr <=  "0001110100001";
		Trees_din <= x"fffe0ec9";
		wait for Clk_period;
		Addr <=  "0001110100010";
		Trees_din <= x"ffcf0ec9";
		wait for Clk_period;
		Addr <=  "0001110100011";
		Trees_din <= x"0cfed404";
		wait for Clk_period;
		Addr <=  "0001110100100";
		Trees_din <= x"ff740ec9";
		wait for Clk_period;
		Addr <=  "0001110100101";
		Trees_din <= x"34ffd610";
		wait for Clk_period;
		Addr <=  "0001110100110";
		Trees_din <= x"57ff4d08";
		wait for Clk_period;
		Addr <=  "0001110100111";
		Trees_din <= x"ccffb004";
		wait for Clk_period;
		Addr <=  "0001110101000";
		Trees_din <= x"00800ec9";
		wait for Clk_period;
		Addr <=  "0001110101001";
		Trees_din <= x"ffd30ec9";
		wait for Clk_period;
		Addr <=  "0001110101010";
		Trees_din <= x"5cffb304";
		wait for Clk_period;
		Addr <=  "0001110101011";
		Trees_din <= x"fff70ec9";
		wait for Clk_period;
		Addr <=  "0001110101100";
		Trees_din <= x"ff930ec9";
		wait for Clk_period;
		Addr <=  "0001110101101";
		Trees_din <= x"4bff7908";
		wait for Clk_period;
		Addr <=  "0001110101110";
		Trees_din <= x"fdff0004";
		wait for Clk_period;
		Addr <=  "0001110101111";
		Trees_din <= x"fffd0ec9";
		wait for Clk_period;
		Addr <=  "0001110110000";
		Trees_din <= x"ff7b0ec9";
		wait for Clk_period;
		Addr <=  "0001110110001";
		Trees_din <= x"00100ec9";
		wait for Clk_period;
		Addr <=  "0001110110010";
		Trees_din <= x"14ff4a14";
		wait for Clk_period;
		Addr <=  "0001110110011";
		Trees_din <= x"9dfeb308";
		wait for Clk_period;
		Addr <=  "0001110110100";
		Trees_din <= x"e1003b04";
		wait for Clk_period;
		Addr <=  "0001110110101";
		Trees_din <= x"ffb00f65";
		wait for Clk_period;
		Addr <=  "0001110110110";
		Trees_din <= x"007d0f65";
		wait for Clk_period;
		Addr <=  "0001110110111";
		Trees_din <= x"d2ff5804";
		wait for Clk_period;
		Addr <=  "0001110111000";
		Trees_din <= x"ff690f65";
		wait for Clk_period;
		Addr <=  "0001110111001";
		Trees_din <= x"fe001b04";
		wait for Clk_period;
		Addr <=  "0001110111010";
		Trees_din <= x"ff960f65";
		wait for Clk_period;
		Addr <=  "0001110111011";
		Trees_din <= x"00360f65";
		wait for Clk_period;
		Addr <=  "0001110111100";
		Trees_din <= x"13004f24";
		wait for Clk_period;
		Addr <=  "0001110111101";
		Trees_din <= x"e2ff8e1c";
		wait for Clk_period;
		Addr <=  "0001110111110";
		Trees_din <= x"83ff520c";
		wait for Clk_period;
		Addr <=  "0001110111111";
		Trees_din <= x"bd007c08";
		wait for Clk_period;
		Addr <=  "0001111000000";
		Trees_din <= x"76ffc804";
		wait for Clk_period;
		Addr <=  "0001111000001";
		Trees_din <= x"00160f65";
		wait for Clk_period;
		Addr <=  "0001111000010";
		Trees_din <= x"00990f65";
		wait for Clk_period;
		Addr <=  "0001111000011";
		Trees_din <= x"ffdf0f65";
		wait for Clk_period;
		Addr <=  "0001111000100";
		Trees_din <= x"eafff108";
		wait for Clk_period;
		Addr <=  "0001111000101";
		Trees_din <= x"f7feed04";
		wait for Clk_period;
		Addr <=  "0001111000110";
		Trees_din <= x"00330f65";
		wait for Clk_period;
		Addr <=  "0001111000111";
		Trees_din <= x"ff9b0f65";
		wait for Clk_period;
		Addr <=  "0001111001000";
		Trees_din <= x"7fff8204";
		wait for Clk_period;
		Addr <=  "0001111001001";
		Trees_din <= x"005b0f65";
		wait for Clk_period;
		Addr <=  "0001111001010";
		Trees_din <= x"000e0f65";
		wait for Clk_period;
		Addr <=  "0001111001011";
		Trees_din <= x"e3ff3904";
		wait for Clk_period;
		Addr <=  "0001111001100";
		Trees_din <= x"ff8b0f65";
		wait for Clk_period;
		Addr <=  "0001111001101";
		Trees_din <= x"004b0f65";
		wait for Clk_period;
		Addr <=  "0001111001110";
		Trees_din <= x"0eff0e08";
		wait for Clk_period;
		Addr <=  "0001111001111";
		Trees_din <= x"ddfeaf04";
		wait for Clk_period;
		Addr <=  "0001111010000";
		Trees_din <= x"fff40f65";
		wait for Clk_period;
		Addr <=  "0001111010001";
		Trees_din <= x"ff770f65";
		wait for Clk_period;
		Addr <=  "0001111010010";
		Trees_din <= x"0cfed404";
		wait for Clk_period;
		Addr <=  "0001111010011";
		Trees_din <= x"ff8d0f65";
		wait for Clk_period;
		Addr <=  "0001111010100";
		Trees_din <= x"31ffad08";
		wait for Clk_period;
		Addr <=  "0001111010101";
		Trees_din <= x"d9ffe504";
		wait for Clk_period;
		Addr <=  "0001111010110";
		Trees_din <= x"006d0f65";
		wait for Clk_period;
		Addr <=  "0001111010111";
		Trees_din <= x"ffdb0f65";
		wait for Clk_period;
		Addr <=  "0001111011000";
		Trees_din <= x"ffa90f65";
		wait for Clk_period;
		Addr <=  "0001111011001";
		Trees_din <= x"14ff4a10";
		wait for Clk_period;
		Addr <=  "0001111011010";
		Trees_din <= x"9dfeb304";
		wait for Clk_period;
		Addr <=  "0001111011011";
		Trees_din <= x"001d1031";
		wait for Clk_period;
		Addr <=  "0001111011100";
		Trees_din <= x"d2ff5804";
		wait for Clk_period;
		Addr <=  "0001111011101";
		Trees_din <= x"ff6a1031";
		wait for Clk_period;
		Addr <=  "0001111011110";
		Trees_din <= x"e8001f04";
		wait for Clk_period;
		Addr <=  "0001111011111";
		Trees_din <= x"ff9a1031";
		wait for Clk_period;
		Addr <=  "0001111100000";
		Trees_din <= x"00341031";
		wait for Clk_period;
		Addr <=  "0001111100001";
		Trees_din <= x"13004f30";
		wait for Clk_period;
		Addr <=  "0001111100010";
		Trees_din <= x"85fff314";
		wait for Clk_period;
		Addr <=  "0001111100011";
		Trees_din <= x"1700450c";
		wait for Clk_period;
		Addr <=  "0001111100100";
		Trees_din <= x"7500a308";
		wait for Clk_period;
		Addr <=  "0001111100101";
		Trees_din <= x"b7ff8004";
		wait for Clk_period;
		Addr <=  "0001111100110";
		Trees_din <= x"000d1031";
		wait for Clk_period;
		Addr <=  "0001111100111";
		Trees_din <= x"ff881031";
		wait for Clk_period;
		Addr <=  "0001111101000";
		Trees_din <= x"004b1031";
		wait for Clk_period;
		Addr <=  "0001111101001";
		Trees_din <= x"78ffae04";
		wait for Clk_period;
		Addr <=  "0001111101010";
		Trees_din <= x"ffff1031";
		wait for Clk_period;
		Addr <=  "0001111101011";
		Trees_din <= x"007e1031";
		wait for Clk_period;
		Addr <=  "0001111101100";
		Trees_din <= x"03ff630c";
		wait for Clk_period;
		Addr <=  "0001111101101";
		Trees_din <= x"96ff6b04";
		wait for Clk_period;
		Addr <=  "0001111101110";
		Trees_din <= x"001c1031";
		wait for Clk_period;
		Addr <=  "0001111101111";
		Trees_din <= x"26001b04";
		wait for Clk_period;
		Addr <=  "0001111110000";
		Trees_din <= x"002e1031";
		wait for Clk_period;
		Addr <=  "0001111110001";
		Trees_din <= x"00a11031";
		wait for Clk_period;
		Addr <=  "0001111110010";
		Trees_din <= x"29001c08";
		wait for Clk_period;
		Addr <=  "0001111110011";
		Trees_din <= x"52feef04";
		wait for Clk_period;
		Addr <=  "0001111110100";
		Trees_din <= x"00251031";
		wait for Clk_period;
		Addr <=  "0001111110101";
		Trees_din <= x"ff9d1031";
		wait for Clk_period;
		Addr <=  "0001111110110";
		Trees_din <= x"b0ffed04";
		wait for Clk_period;
		Addr <=  "0001111110111";
		Trees_din <= x"006f1031";
		wait for Clk_period;
		Addr <=  "0001111111000";
		Trees_din <= x"fffe1031";
		wait for Clk_period;
		Addr <=  "0001111111001";
		Trees_din <= x"0eff5c14";
		wait for Clk_period;
		Addr <=  "0001111111010";
		Trees_din <= x"4f002908";
		wait for Clk_period;
		Addr <=  "0001111111011";
		Trees_din <= x"5e003b04";
		wait for Clk_period;
		Addr <=  "0001111111100";
		Trees_din <= x"ff781031";
		wait for Clk_period;
		Addr <=  "0001111111101";
		Trees_din <= x"ffed1031";
		wait for Clk_period;
		Addr <=  "0001111111110";
		Trees_din <= x"a0ff6804";
		wait for Clk_period;
		Addr <=  "0001111111111";
		Trees_din <= x"ffa71031";
		wait for Clk_period;
		Addr <=  "0010000000000";
		Trees_din <= x"e3fed504";
		wait for Clk_period;
		Addr <=  "0010000000001";
		Trees_din <= x"ffed1031";
		wait for Clk_period;
		Addr <=  "0010000000010";
		Trees_din <= x"00631031";
		wait for Clk_period;
		Addr <=  "0010000000011";
		Trees_din <= x"70ff5008";
		wait for Clk_period;
		Addr <=  "0010000000100";
		Trees_din <= x"88000304";
		wait for Clk_period;
		Addr <=  "0010000000101";
		Trees_din <= x"ffa51031";
		wait for Clk_period;
		Addr <=  "0010000000110";
		Trees_din <= x"ffeb1031";
		wait for Clk_period;
		Addr <=  "0010000000111";
		Trees_din <= x"6affd408";
		wait for Clk_period;
		Addr <=  "0010000001000";
		Trees_din <= x"c2ff2704";
		wait for Clk_period;
		Addr <=  "0010000001001";
		Trees_din <= x"00931031";
		wait for Clk_period;
		Addr <=  "0010000001010";
		Trees_din <= x"00281031";
		wait for Clk_period;
		Addr <=  "0010000001011";
		Trees_din <= x"ffd11031";
		wait for Clk_period;
		Addr <=  "0010000001100";
		Trees_din <= x"0eff0e18";
		wait for Clk_period;
		Addr <=  "0010000001101";
		Trees_din <= x"0cffc20c";
		wait for Clk_period;
		Addr <=  "0010000001110";
		Trees_din <= x"92fff708";
		wait for Clk_period;
		Addr <=  "0010000001111";
		Trees_din <= x"aefe0004";
		wait for Clk_period;
		Addr <=  "0010000010000";
		Trees_din <= x"ffe910c5";
		wait for Clk_period;
		Addr <=  "0010000010001";
		Trees_din <= x"ff6a10c5";
		wait for Clk_period;
		Addr <=  "0010000010010";
		Trees_din <= x"001a10c5";
		wait for Clk_period;
		Addr <=  "0010000010011";
		Trees_din <= x"85ffd504";
		wait for Clk_period;
		Addr <=  "0010000010100";
		Trees_din <= x"ffab10c5";
		wait for Clk_period;
		Addr <=  "0010000010101";
		Trees_din <= x"b7ffc904";
		wait for Clk_period;
		Addr <=  "0010000010110";
		Trees_din <= x"ffff10c5";
		wait for Clk_period;
		Addr <=  "0010000010111";
		Trees_din <= x"007110c5";
		wait for Clk_period;
		Addr <=  "0010000011000";
		Trees_din <= x"baff9714";
		wait for Clk_period;
		Addr <=  "0010000011001";
		Trees_din <= x"92ff1b04";
		wait for Clk_period;
		Addr <=  "0010000011010";
		Trees_din <= x"ff9c10c5";
		wait for Clk_period;
		Addr <=  "0010000011011";
		Trees_din <= x"57ff970c";
		wait for Clk_period;
		Addr <=  "0010000011100";
		Trees_din <= x"4eff4204";
		wait for Clk_period;
		Addr <=  "0010000011101";
		Trees_din <= x"ffcb10c5";
		wait for Clk_period;
		Addr <=  "0010000011110";
		Trees_din <= x"b2001304";
		wait for Clk_period;
		Addr <=  "0010000011111";
		Trees_din <= x"008d10c5";
		wait for Clk_period;
		Addr <=  "0010000100000";
		Trees_din <= x"fffe10c5";
		wait for Clk_period;
		Addr <=  "0010000100001";
		Trees_din <= x"ffc810c5";
		wait for Clk_period;
		Addr <=  "0010000100010";
		Trees_din <= x"76001210";
		wait for Clk_period;
		Addr <=  "0010000100011";
		Trees_din <= x"e8003f08";
		wait for Clk_period;
		Addr <=  "0010000100100";
		Trees_din <= x"36ffc604";
		wait for Clk_period;
		Addr <=  "0010000100101";
		Trees_din <= x"ff7810c5";
		wait for Clk_period;
		Addr <=  "0010000100110";
		Trees_din <= x"ffe410c5";
		wait for Clk_period;
		Addr <=  "0010000100111";
		Trees_din <= x"5dffb204";
		wait for Clk_period;
		Addr <=  "0010000101000";
		Trees_din <= x"ffb110c5";
		wait for Clk_period;
		Addr <=  "0010000101001";
		Trees_din <= x"003c10c5";
		wait for Clk_period;
		Addr <=  "0010000101010";
		Trees_din <= x"f1ff9e04";
		wait for Clk_period;
		Addr <=  "0010000101011";
		Trees_din <= x"ffad10c5";
		wait for Clk_period;
		Addr <=  "0010000101100";
		Trees_din <= x"8efff708";
		wait for Clk_period;
		Addr <=  "0010000101101";
		Trees_din <= x"70ff2f04";
		wait for Clk_period;
		Addr <=  "0010000101110";
		Trees_din <= x"001b10c5";
		wait for Clk_period;
		Addr <=  "0010000101111";
		Trees_din <= x"007d10c5";
		wait for Clk_period;
		Addr <=  "0010000110000";
		Trees_din <= x"ffd610c5";
		wait for Clk_period;
		Addr <=  "0010000110001";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0010000110010";
		Trees_din <= x"0eff0e14";
		wait for Clk_period;
		Addr <=  "0010000110011";
		Trees_din <= x"0cffc20c";
		wait for Clk_period;
		Addr <=  "0010000110100";
		Trees_din <= x"92fff708";
		wait for Clk_period;
		Addr <=  "0010000110101";
		Trees_din <= x"aefe0004";
		wait for Clk_period;
		Addr <=  "0010000110110";
		Trees_din <= x"ffea114d";
		wait for Clk_period;
		Addr <=  "0010000110111";
		Trees_din <= x"ff6b114d";
		wait for Clk_period;
		Addr <=  "0010000111000";
		Trees_din <= x"0016114d";
		wait for Clk_period;
		Addr <=  "0010000111001";
		Trees_din <= x"e3ff1404";
		wait for Clk_period;
		Addr <=  "0010000111010";
		Trees_din <= x"ffbf114d";
		wait for Clk_period;
		Addr <=  "0010000111011";
		Trees_din <= x"005b114d";
		wait for Clk_period;
		Addr <=  "0010000111100";
		Trees_din <= x"b0ff6f08";
		wait for Clk_period;
		Addr <=  "0010000111101";
		Trees_din <= x"8cff1a04";
		wait for Clk_period;
		Addr <=  "0010000111110";
		Trees_din <= x"0003114d";
		wait for Clk_period;
		Addr <=  "0010000111111";
		Trees_din <= x"ff80114d";
		wait for Clk_period;
		Addr <=  "0010001000000";
		Trees_din <= x"1300d520";
		wait for Clk_period;
		Addr <=  "0010001000001";
		Trees_din <= x"baff9710";
		wait for Clk_period;
		Addr <=  "0010001000010";
		Trees_din <= x"e2ff7608";
		wait for Clk_period;
		Addr <=  "0010001000011";
		Trees_din <= x"b2001304";
		wait for Clk_period;
		Addr <=  "0010001000100";
		Trees_din <= x"0090114d";
		wait for Clk_period;
		Addr <=  "0010001000101";
		Trees_din <= x"fff0114d";
		wait for Clk_period;
		Addr <=  "0010001000110";
		Trees_din <= x"6cff3a04";
		wait for Clk_period;
		Addr <=  "0010001000111";
		Trees_din <= x"003e114d";
		wait for Clk_period;
		Addr <=  "0010001001000";
		Trees_din <= x"ffc0114d";
		wait for Clk_period;
		Addr <=  "0010001001001";
		Trees_din <= x"c2ff3f08";
		wait for Clk_period;
		Addr <=  "0010001001010";
		Trees_din <= x"34ffd804";
		wait for Clk_period;
		Addr <=  "0010001001011";
		Trees_din <= x"0056114d";
		wait for Clk_period;
		Addr <=  "0010001001100";
		Trees_din <= x"ffdc114d";
		wait for Clk_period;
		Addr <=  "0010001001101";
		Trees_din <= x"3fffe704";
		wait for Clk_period;
		Addr <=  "0010001001110";
		Trees_din <= x"0014114d";
		wait for Clk_period;
		Addr <=  "0010001001111";
		Trees_din <= x"ff93114d";
		wait for Clk_period;
		Addr <=  "0010001010000";
		Trees_din <= x"a3ff2604";
		wait for Clk_period;
		Addr <=  "0010001010001";
		Trees_din <= x"fffc114d";
		wait for Clk_period;
		Addr <=  "0010001010010";
		Trees_din <= x"ff92114d";
		wait for Clk_period;
		Addr <=  "0010001010011";
		Trees_din <= x"70ff2418";
		wait for Clk_period;
		Addr <=  "0010001010100";
		Trees_din <= x"ebff6008";
		wait for Clk_period;
		Addr <=  "0010001010101";
		Trees_din <= x"95001504";
		wait for Clk_period;
		Addr <=  "0010001010110";
		Trees_din <= x"ff6c11e9";
		wait for Clk_period;
		Addr <=  "0010001010111";
		Trees_din <= x"001b11e9";
		wait for Clk_period;
		Addr <=  "0010001011000";
		Trees_din <= x"84005608";
		wait for Clk_period;
		Addr <=  "0010001011001";
		Trees_din <= x"f1000f04";
		wait for Clk_period;
		Addr <=  "0010001011010";
		Trees_din <= x"ff9b11e9";
		wait for Clk_period;
		Addr <=  "0010001011011";
		Trees_din <= x"001211e9";
		wait for Clk_period;
		Addr <=  "0010001011100";
		Trees_din <= x"5cffd404";
		wait for Clk_period;
		Addr <=  "0010001011101";
		Trees_din <= x"007211e9";
		wait for Clk_period;
		Addr <=  "0010001011110";
		Trees_din <= x"001711e9";
		wait for Clk_period;
		Addr <=  "0010001011111";
		Trees_din <= x"34ffd620";
		wait for Clk_period;
		Addr <=  "0010001100000";
		Trees_din <= x"15ff4008";
		wait for Clk_period;
		Addr <=  "0010001100001";
		Trees_din <= x"51002004";
		wait for Clk_period;
		Addr <=  "0010001100010";
		Trees_din <= x"ff9a11e9";
		wait for Clk_period;
		Addr <=  "0010001100011";
		Trees_din <= x"002d11e9";
		wait for Clk_period;
		Addr <=  "0010001100100";
		Trees_din <= x"72ffbf08";
		wait for Clk_period;
		Addr <=  "0010001100101";
		Trees_din <= x"c1ff1704";
		wait for Clk_period;
		Addr <=  "0010001100110";
		Trees_din <= x"ffa611e9";
		wait for Clk_period;
		Addr <=  "0010001100111";
		Trees_din <= x"001a11e9";
		wait for Clk_period;
		Addr <=  "0010001101000";
		Trees_din <= x"c2ff7808";
		wait for Clk_period;
		Addr <=  "0010001101001";
		Trees_din <= x"f1ff8c04";
		wait for Clk_period;
		Addr <=  "0010001101010";
		Trees_din <= x"001011e9";
		wait for Clk_period;
		Addr <=  "0010001101011";
		Trees_din <= x"009411e9";
		wait for Clk_period;
		Addr <=  "0010001101100";
		Trees_din <= x"d2ff3704";
		wait for Clk_period;
		Addr <=  "0010001101101";
		Trees_din <= x"ffcd11e9";
		wait for Clk_period;
		Addr <=  "0010001101110";
		Trees_din <= x"003b11e9";
		wait for Clk_period;
		Addr <=  "0010001101111";
		Trees_din <= x"ebff6308";
		wait for Clk_period;
		Addr <=  "0010001110000";
		Trees_din <= x"13001b04";
		wait for Clk_period;
		Addr <=  "0010001110001";
		Trees_din <= x"fffb11e9";
		wait for Clk_period;
		Addr <=  "0010001110010";
		Trees_din <= x"ff7a11e9";
		wait for Clk_period;
		Addr <=  "0010001110011";
		Trees_din <= x"baff9708";
		wait for Clk_period;
		Addr <=  "0010001110100";
		Trees_din <= x"f7ff6a04";
		wait for Clk_period;
		Addr <=  "0010001110101";
		Trees_din <= x"007611e9";
		wait for Clk_period;
		Addr <=  "0010001110110";
		Trees_din <= x"fff511e9";
		wait for Clk_period;
		Addr <=  "0010001110111";
		Trees_din <= x"b9ff3c04";
		wait for Clk_period;
		Addr <=  "0010001111000";
		Trees_din <= x"000c11e9";
		wait for Clk_period;
		Addr <=  "0010001111001";
		Trees_din <= x"ffaf11e9";
		wait for Clk_period;
		Addr <=  "0010001111010";
		Trees_din <= x"14ff480c";
		wait for Clk_period;
		Addr <=  "0010001111011";
		Trees_din <= x"9dfeb304";
		wait for Clk_period;
		Addr <=  "0010001111100";
		Trees_din <= x"0021127d";
		wait for Clk_period;
		Addr <=  "0010001111101";
		Trees_din <= x"e3ff4404";
		wait for Clk_period;
		Addr <=  "0010001111110";
		Trees_din <= x"ff6e127d";
		wait for Clk_period;
		Addr <=  "0010001111111";
		Trees_din <= x"fff2127d";
		wait for Clk_period;
		Addr <=  "0010010000000";
		Trees_din <= x"13004f24";
		wait for Clk_period;
		Addr <=  "0010010000001";
		Trees_din <= x"96ffc410";
		wait for Clk_period;
		Addr <=  "0010010000010";
		Trees_din <= x"e9ff8308";
		wait for Clk_period;
		Addr <=  "0010010000011";
		Trees_din <= x"c6ffc804";
		wait for Clk_period;
		Addr <=  "0010010000100";
		Trees_din <= x"ff9a127d";
		wait for Clk_period;
		Addr <=  "0010010000101";
		Trees_din <= x"002c127d";
		wait for Clk_period;
		Addr <=  "0010010000110";
		Trees_din <= x"b2ff9e04";
		wait for Clk_period;
		Addr <=  "0010010000111";
		Trees_din <= x"ffed127d";
		wait for Clk_period;
		Addr <=  "0010010001000";
		Trees_din <= x"0062127d";
		wait for Clk_period;
		Addr <=  "0010010001001";
		Trees_din <= x"78ff7308";
		wait for Clk_period;
		Addr <=  "0010010001010";
		Trees_din <= x"74ffd304";
		wait for Clk_period;
		Addr <=  "0010010001011";
		Trees_din <= x"ffbb127d";
		wait for Clk_period;
		Addr <=  "0010010001100";
		Trees_din <= x"0028127d";
		wait for Clk_period;
		Addr <=  "0010010001101";
		Trees_din <= x"83ff6608";
		wait for Clk_period;
		Addr <=  "0010010001110";
		Trees_din <= x"25003204";
		wait for Clk_period;
		Addr <=  "0010010001111";
		Trees_din <= x"009a127d";
		wait for Clk_period;
		Addr <=  "0010010010000";
		Trees_din <= x"0030127d";
		wait for Clk_period;
		Addr <=  "0010010010001";
		Trees_din <= x"0005127d";
		wait for Clk_period;
		Addr <=  "0010010010010";
		Trees_din <= x"0cfed404";
		wait for Clk_period;
		Addr <=  "0010010010011";
		Trees_din <= x"ff84127d";
		wait for Clk_period;
		Addr <=  "0010010010100";
		Trees_din <= x"b8002910";
		wait for Clk_period;
		Addr <=  "0010010010101";
		Trees_din <= x"dfffb808";
		wait for Clk_period;
		Addr <=  "0010010010110";
		Trees_din <= x"86ffda04";
		wait for Clk_period;
		Addr <=  "0010010010111";
		Trees_din <= x"ff86127d";
		wait for Clk_period;
		Addr <=  "0010010011000";
		Trees_din <= x"002a127d";
		wait for Clk_period;
		Addr <=  "0010010011001";
		Trees_din <= x"c5ff7104";
		wait for Clk_period;
		Addr <=  "0010010011010";
		Trees_din <= x"fffe127d";
		wait for Clk_period;
		Addr <=  "0010010011011";
		Trees_din <= x"0050127d";
		wait for Clk_period;
		Addr <=  "0010010011100";
		Trees_din <= x"baff7a04";
		wait for Clk_period;
		Addr <=  "0010010011101";
		Trees_din <= x"006d127d";
		wait for Clk_period;
		Addr <=  "0010010011110";
		Trees_din <= x"fffd127d";
		wait for Clk_period;
		Addr <=  "0010010011111";
		Trees_din <= x"70ff2414";
		wait for Clk_period;
		Addr <=  "0010010100000";
		Trees_din <= x"ebff6008";
		wait for Clk_period;
		Addr <=  "0010010100001";
		Trees_din <= x"a5fe8a04";
		wait for Clk_period;
		Addr <=  "0010010100010";
		Trees_din <= x"00011301";
		wait for Clk_period;
		Addr <=  "0010010100011";
		Trees_din <= x"ff701301";
		wait for Clk_period;
		Addr <=  "0010010100100";
		Trees_din <= x"84005608";
		wait for Clk_period;
		Addr <=  "0010010100101";
		Trees_din <= x"f1fffc04";
		wait for Clk_period;
		Addr <=  "0010010100110";
		Trees_din <= x"ffa11301";
		wait for Clk_period;
		Addr <=  "0010010100111";
		Trees_din <= x"000f1301";
		wait for Clk_period;
		Addr <=  "0010010101000";
		Trees_din <= x"00511301";
		wait for Clk_period;
		Addr <=  "0010010101001";
		Trees_din <= x"85fff51c";
		wait for Clk_period;
		Addr <=  "0010010101010";
		Trees_din <= x"92ffd610";
		wait for Clk_period;
		Addr <=  "0010010101011";
		Trees_din <= x"baff6508";
		wait for Clk_period;
		Addr <=  "0010010101100";
		Trees_din <= x"0eff6104";
		wait for Clk_period;
		Addr <=  "0010010101101";
		Trees_din <= x"ffc71301";
		wait for Clk_period;
		Addr <=  "0010010101110";
		Trees_din <= x"00461301";
		wait for Clk_period;
		Addr <=  "0010010101111";
		Trees_din <= x"96ffee04";
		wait for Clk_period;
		Addr <=  "0010010110000";
		Trees_din <= x"ff7d1301";
		wait for Clk_period;
		Addr <=  "0010010110001";
		Trees_din <= x"ffe21301";
		wait for Clk_period;
		Addr <=  "0010010110010";
		Trees_din <= x"f1ffa904";
		wait for Clk_period;
		Addr <=  "0010010110011";
		Trees_din <= x"ffcd1301";
		wait for Clk_period;
		Addr <=  "0010010110100";
		Trees_din <= x"27ffc104";
		wait for Clk_period;
		Addr <=  "0010010110101";
		Trees_din <= x"001b1301";
		wait for Clk_period;
		Addr <=  "0010010110110";
		Trees_din <= x"00771301";
		wait for Clk_period;
		Addr <=  "0010010110111";
		Trees_din <= x"15ff3804";
		wait for Clk_period;
		Addr <=  "0010010111000";
		Trees_din <= x"ffb61301";
		wait for Clk_period;
		Addr <=  "0010010111001";
		Trees_din <= x"83ff950c";
		wait for Clk_period;
		Addr <=  "0010010111010";
		Trees_din <= x"f9ff6208";
		wait for Clk_period;
		Addr <=  "0010010111011";
		Trees_din <= x"bcfefc04";
		wait for Clk_period;
		Addr <=  "0010010111100";
		Trees_din <= x"000d1301";
		wait for Clk_period;
		Addr <=  "0010010111101";
		Trees_din <= x"008e1301";
		wait for Clk_period;
		Addr <=  "0010010111110";
		Trees_din <= x"fff51301";
		wait for Clk_period;
		Addr <=  "0010010111111";
		Trees_din <= x"ffdb1301";
		wait for Clk_period;
		Addr <=  "0010011000000";
		Trees_din <= x"0eff0014";
		wait for Clk_period;
		Addr <=  "0010011000001";
		Trees_din <= x"0cffc20c";
		wait for Clk_period;
		Addr <=  "0010011000010";
		Trees_din <= x"92fff708";
		wait for Clk_period;
		Addr <=  "0010011000011";
		Trees_din <= x"d800a704";
		wait for Clk_period;
		Addr <=  "0010011000100";
		Trees_din <= x"ff70137d";
		wait for Clk_period;
		Addr <=  "0010011000101";
		Trees_din <= x"ffdb137d";
		wait for Clk_period;
		Addr <=  "0010011000110";
		Trees_din <= x"0009137d";
		wait for Clk_period;
		Addr <=  "0010011000111";
		Trees_din <= x"e3ff1404";
		wait for Clk_period;
		Addr <=  "0010011001000";
		Trees_din <= x"ffd4137d";
		wait for Clk_period;
		Addr <=  "0010011001001";
		Trees_din <= x"0041137d";
		wait for Clk_period;
		Addr <=  "0010011001010";
		Trees_din <= x"70ff100c";
		wait for Clk_period;
		Addr <=  "0010011001011";
		Trees_din <= x"84008a08";
		wait for Clk_period;
		Addr <=  "0010011001100";
		Trees_din <= x"11000f04";
		wait for Clk_period;
		Addr <=  "0010011001101";
		Trees_din <= x"ff85137d";
		wait for Clk_period;
		Addr <=  "0010011001110";
		Trees_din <= x"0010137d";
		wait for Clk_period;
		Addr <=  "0010011001111";
		Trees_din <= x"003c137d";
		wait for Clk_period;
		Addr <=  "0010011010000";
		Trees_din <= x"baff9710";
		wait for Clk_period;
		Addr <=  "0010011010001";
		Trees_din <= x"15ff3804";
		wait for Clk_period;
		Addr <=  "0010011010010";
		Trees_din <= x"ffdd137d";
		wait for Clk_period;
		Addr <=  "0010011010011";
		Trees_din <= x"e5fe8c04";
		wait for Clk_period;
		Addr <=  "0010011010100";
		Trees_din <= x"fff5137d";
		wait for Clk_period;
		Addr <=  "0010011010101";
		Trees_din <= x"8b000104";
		wait for Clk_period;
		Addr <=  "0010011010110";
		Trees_din <= x"008b137d";
		wait for Clk_period;
		Addr <=  "0010011010111";
		Trees_din <= x"0016137d";
		wait for Clk_period;
		Addr <=  "0010011011000";
		Trees_din <= x"97fef808";
		wait for Clk_period;
		Addr <=  "0010011011001";
		Trees_din <= x"cbfff104";
		wait for Clk_period;
		Addr <=  "0010011011010";
		Trees_din <= x"fff0137d";
		wait for Clk_period;
		Addr <=  "0010011011011";
		Trees_din <= x"0057137d";
		wait for Clk_period;
		Addr <=  "0010011011100";
		Trees_din <= x"76002704";
		wait for Clk_period;
		Addr <=  "0010011011101";
		Trees_din <= x"ff9a137d";
		wait for Clk_period;
		Addr <=  "0010011011110";
		Trees_din <= x"000e137d";
		wait for Clk_period;
		Addr <=  "0010011011111";
		Trees_din <= x"0eff0014";
		wait for Clk_period;
		Addr <=  "0010011100000";
		Trees_din <= x"34ffb90c";
		wait for Clk_period;
		Addr <=  "0010011100001";
		Trees_din <= x"c0ffa604";
		wait for Clk_period;
		Addr <=  "0010011100010";
		Trees_din <= x"ffb313f1";
		wait for Clk_period;
		Addr <=  "0010011100011";
		Trees_din <= x"a7ff9d04";
		wait for Clk_period;
		Addr <=  "0010011100100";
		Trees_din <= x"004f13f1";
		wait for Clk_period;
		Addr <=  "0010011100101";
		Trees_din <= x"fffb13f1";
		wait for Clk_period;
		Addr <=  "0010011100110";
		Trees_din <= x"84004804";
		wait for Clk_period;
		Addr <=  "0010011100111";
		Trees_din <= x"ff7313f1";
		wait for Clk_period;
		Addr <=  "0010011101000";
		Trees_din <= x"ffd113f1";
		wait for Clk_period;
		Addr <=  "0010011101001";
		Trees_din <= x"1300d520";
		wait for Clk_period;
		Addr <=  "0010011101010";
		Trees_din <= x"bcfefc08";
		wait for Clk_period;
		Addr <=  "0010011101011";
		Trees_din <= x"92fff104";
		wait for Clk_period;
		Addr <=  "0010011101100";
		Trees_din <= x"ffa613f1";
		wait for Clk_period;
		Addr <=  "0010011101101";
		Trees_din <= x"001f13f1";
		wait for Clk_period;
		Addr <=  "0010011101110";
		Trees_din <= x"e2ff740c";
		wait for Clk_period;
		Addr <=  "0010011101111";
		Trees_din <= x"bd006a08";
		wait for Clk_period;
		Addr <=  "0010011110000";
		Trees_din <= x"b2001304";
		wait for Clk_period;
		Addr <=  "0010011110001";
		Trees_din <= x"006d13f1";
		wait for Clk_period;
		Addr <=  "0010011110010";
		Trees_din <= x"ffea13f1";
		wait for Clk_period;
		Addr <=  "0010011110011";
		Trees_din <= x"ffcb13f1";
		wait for Clk_period;
		Addr <=  "0010011110100";
		Trees_din <= x"51002808";
		wait for Clk_period;
		Addr <=  "0010011110101";
		Trees_din <= x"adff9804";
		wait for Clk_period;
		Addr <=  "0010011110110";
		Trees_din <= x"ffa813f1";
		wait for Clk_period;
		Addr <=  "0010011110111";
		Trees_din <= x"001213f1";
		wait for Clk_period;
		Addr <=  "0010011111000";
		Trees_din <= x"004613f1";
		wait for Clk_period;
		Addr <=  "0010011111001";
		Trees_din <= x"c5ff8904";
		wait for Clk_period;
		Addr <=  "0010011111010";
		Trees_din <= x"ff9113f1";
		wait for Clk_period;
		Addr <=  "0010011111011";
		Trees_din <= x"000913f1";
		wait for Clk_period;
		Addr <=  "0010011111100";
		Trees_din <= x"70ff2410";
		wait for Clk_period;
		Addr <=  "0010011111101";
		Trees_din <= x"ebff6008";
		wait for Clk_period;
		Addr <=  "0010011111110";
		Trees_din <= x"6bff3d04";
		wait for Clk_period;
		Addr <=  "0010011111111";
		Trees_din <= x"ff761465";
		wait for Clk_period;
		Addr <=  "0010100000000";
		Trees_din <= x"ffd81465";
		wait for Clk_period;
		Addr <=  "0010100000001";
		Trees_din <= x"d2ff4f04";
		wait for Clk_period;
		Addr <=  "0010100000010";
		Trees_din <= x"ffcb1465";
		wait for Clk_period;
		Addr <=  "0010100000011";
		Trees_din <= x"00491465";
		wait for Clk_period;
		Addr <=  "0010100000100";
		Trees_din <= x"85fff514";
		wait for Clk_period;
		Addr <=  "0010100000101";
		Trees_din <= x"92ffd60c";
		wait for Clk_period;
		Addr <=  "0010100000110";
		Trees_din <= x"baff6504";
		wait for Clk_period;
		Addr <=  "0010100000111";
		Trees_din <= x"000d1465";
		wait for Clk_period;
		Addr <=  "0010100001000";
		Trees_din <= x"96ffee04";
		wait for Clk_period;
		Addr <=  "0010100001001";
		Trees_din <= x"ff861465";
		wait for Clk_period;
		Addr <=  "0010100001010";
		Trees_din <= x"ffe61465";
		wait for Clk_period;
		Addr <=  "0010100001011";
		Trees_din <= x"d2ff1604";
		wait for Clk_period;
		Addr <=  "0010100001100";
		Trees_din <= x"00581465";
		wait for Clk_period;
		Addr <=  "0010100001101";
		Trees_din <= x"ffd81465";
		wait for Clk_period;
		Addr <=  "0010100001110";
		Trees_din <= x"03ff830c";
		wait for Clk_period;
		Addr <=  "0010100001111";
		Trees_din <= x"fcff5b04";
		wait for Clk_period;
		Addr <=  "0010100010000";
		Trees_din <= x"000a1465";
		wait for Clk_period;
		Addr <=  "0010100010001";
		Trees_din <= x"52ff4304";
		wait for Clk_period;
		Addr <=  "0010100010010";
		Trees_din <= x"00801465";
		wait for Clk_period;
		Addr <=  "0010100010011";
		Trees_din <= x"001b1465";
		wait for Clk_period;
		Addr <=  "0010100010100";
		Trees_din <= x"07ffef04";
		wait for Clk_period;
		Addr <=  "0010100010101";
		Trees_din <= x"003b1465";
		wait for Clk_period;
		Addr <=  "0010100010110";
		Trees_din <= x"4f003504";
		wait for Clk_period;
		Addr <=  "0010100010111";
		Trees_din <= x"ffaf1465";
		wait for Clk_period;
		Addr <=  "0010100011000";
		Trees_din <= x"ffea1465";
		wait for Clk_period;
		Addr <=  "0010100011001";
		Trees_din <= x"13004f20";
		wait for Clk_period;
		Addr <=  "0010100011010";
		Trees_din <= x"ebfee604";
		wait for Clk_period;
		Addr <=  "0010100011011";
		Trees_din <= x"ffbc14d1";
		wait for Clk_period;
		Addr <=  "0010100011100";
		Trees_din <= x"83ff5210";
		wait for Clk_period;
		Addr <=  "0010100011101";
		Trees_din <= x"e2ff910c";
		wait for Clk_period;
		Addr <=  "0010100011110";
		Trees_din <= x"bd005508";
		wait for Clk_period;
		Addr <=  "0010100011111";
		Trees_din <= x"4aff0104";
		wait for Clk_period;
		Addr <=  "0010100100000";
		Trees_din <= x"001614d1";
		wait for Clk_period;
		Addr <=  "0010100100001";
		Trees_din <= x"007814d1";
		wait for Clk_period;
		Addr <=  "0010100100010";
		Trees_din <= x"ffef14d1";
		wait for Clk_period;
		Addr <=  "0010100100011";
		Trees_din <= x"ffe414d1";
		wait for Clk_period;
		Addr <=  "0010100100100";
		Trees_din <= x"5a003e04";
		wait for Clk_period;
		Addr <=  "0010100100101";
		Trees_din <= x"002d14d1";
		wait for Clk_period;
		Addr <=  "0010100100110";
		Trees_din <= x"e7ff8d04";
		wait for Clk_period;
		Addr <=  "0010100100111";
		Trees_din <= x"000514d1";
		wait for Clk_period;
		Addr <=  "0010100101000";
		Trees_din <= x"ffb014d1";
		wait for Clk_period;
		Addr <=  "0010100101001";
		Trees_din <= x"34ffd310";
		wait for Clk_period;
		Addr <=  "0010100101010";
		Trees_din <= x"70ff1e04";
		wait for Clk_period;
		Addr <=  "0010100101011";
		Trees_din <= x"ffa314d1";
		wait for Clk_period;
		Addr <=  "0010100101100";
		Trees_din <= x"57ff2d08";
		wait for Clk_period;
		Addr <=  "0010100101101";
		Trees_din <= x"d0007804";
		wait for Clk_period;
		Addr <=  "0010100101110";
		Trees_din <= x"001214d1";
		wait for Clk_period;
		Addr <=  "0010100101111";
		Trees_din <= x"006a14d1";
		wait for Clk_period;
		Addr <=  "0010100110000";
		Trees_din <= x"ffd014d1";
		wait for Clk_period;
		Addr <=  "0010100110001";
		Trees_din <= x"0cffe904";
		wait for Clk_period;
		Addr <=  "0010100110010";
		Trees_din <= x"ff7a14d1";
		wait for Clk_period;
		Addr <=  "0010100110011";
		Trees_din <= x"000514d1";
		wait for Clk_period;
		Addr <=  "0010100110100";
		Trees_din <= x"34ffe920";
		wait for Clk_period;
		Addr <=  "0010100110101";
		Trees_din <= x"e8ff5b04";
		wait for Clk_period;
		Addr <=  "0010100110110";
		Trees_din <= x"ffa21535";
		wait for Clk_period;
		Addr <=  "0010100110111";
		Trees_din <= x"15ff7d0c";
		wait for Clk_period;
		Addr <=  "0010100111000";
		Trees_din <= x"6cffd808";
		wait for Clk_period;
		Addr <=  "0010100111001";
		Trees_din <= x"e1001a04";
		wait for Clk_period;
		Addr <=  "0010100111010";
		Trees_din <= x"ff971535";
		wait for Clk_period;
		Addr <=  "0010100111011";
		Trees_din <= x"000f1535";
		wait for Clk_period;
		Addr <=  "0010100111100";
		Trees_din <= x"005b1535";
		wait for Clk_period;
		Addr <=  "0010100111101";
		Trees_din <= x"aaffd30c";
		wait for Clk_period;
		Addr <=  "0010100111110";
		Trees_din <= x"edfff108";
		wait for Clk_period;
		Addr <=  "0010100111111";
		Trees_din <= x"70ff1604";
		wait for Clk_period;
		Addr <=  "0010101000000";
		Trees_din <= x"000f1535";
		wait for Clk_period;
		Addr <=  "0010101000001";
		Trees_din <= x"00791535";
		wait for Clk_period;
		Addr <=  "0010101000010";
		Trees_din <= x"ffeb1535";
		wait for Clk_period;
		Addr <=  "0010101000011";
		Trees_din <= x"ffea1535";
		wait for Clk_period;
		Addr <=  "0010101000100";
		Trees_din <= x"ebff6b08";
		wait for Clk_period;
		Addr <=  "0010101000101";
		Trees_din <= x"32ff9704";
		wait for Clk_period;
		Addr <=  "0010101000110";
		Trees_din <= x"ff771535";
		wait for Clk_period;
		Addr <=  "0010101000111";
		Trees_din <= x"ffe81535";
		wait for Clk_period;
		Addr <=  "0010101001000";
		Trees_din <= x"83ff3d08";
		wait for Clk_period;
		Addr <=  "0010101001001";
		Trees_din <= x"87ff2104";
		wait for Clk_period;
		Addr <=  "0010101001010";
		Trees_din <= x"00531535";
		wait for Clk_period;
		Addr <=  "0010101001011";
		Trees_din <= x"00011535";
		wait for Clk_period;
		Addr <=  "0010101001100";
		Trees_din <= x"ffda1535";
		wait for Clk_period;
		Addr <=  "0010101001101";
		Trees_din <= x"0eff000c";
		wait for Clk_period;
		Addr <=  "0010101001110";
		Trees_din <= x"0cffc208";
		wait for Clk_period;
		Addr <=  "0010101001111";
		Trees_din <= x"81ff0e04";
		wait for Clk_period;
		Addr <=  "0010101010000";
		Trees_din <= x"fff215a1";
		wait for Clk_period;
		Addr <=  "0010101010001";
		Trees_din <= x"ff7e15a1";
		wait for Clk_period;
		Addr <=  "0010101010010";
		Trees_din <= x"001715a1";
		wait for Clk_period;
		Addr <=  "0010101010011";
		Trees_din <= x"03ffa320";
		wait for Clk_period;
		Addr <=  "0010101010100";
		Trees_din <= x"baff9710";
		wait for Clk_period;
		Addr <=  "0010101010101";
		Trees_din <= x"49fffd0c";
		wait for Clk_period;
		Addr <=  "0010101010110";
		Trees_din <= x"e5fea604";
		wait for Clk_period;
		Addr <=  "0010101010111";
		Trees_din <= x"000a15a1";
		wait for Clk_period;
		Addr <=  "0010101011000";
		Trees_din <= x"4aff2404";
		wait for Clk_period;
		Addr <=  "0010101011001";
		Trees_din <= x"002515a1";
		wait for Clk_period;
		Addr <=  "0010101011010";
		Trees_din <= x"007a15a1";
		wait for Clk_period;
		Addr <=  "0010101011011";
		Trees_din <= x"fff815a1";
		wait for Clk_period;
		Addr <=  "0010101011100";
		Trees_din <= x"97fef808";
		wait for Clk_period;
		Addr <=  "0010101011101";
		Trees_din <= x"cbfff504";
		wait for Clk_period;
		Addr <=  "0010101011110";
		Trees_din <= x"fff815a1";
		wait for Clk_period;
		Addr <=  "0010101011111";
		Trees_din <= x"004a15a1";
		wait for Clk_period;
		Addr <=  "0010101100000";
		Trees_din <= x"1b000a04";
		wait for Clk_period;
		Addr <=  "0010101100001";
		Trees_din <= x"ffab15a1";
		wait for Clk_period;
		Addr <=  "0010101100010";
		Trees_din <= x"000815a1";
		wait for Clk_period;
		Addr <=  "0010101100011";
		Trees_din <= x"14ffd904";
		wait for Clk_period;
		Addr <=  "0010101100100";
		Trees_din <= x"ffa115a1";
		wait for Clk_period;
		Addr <=  "0010101100101";
		Trees_din <= x"36ff3b04";
		wait for Clk_period;
		Addr <=  "0010101100110";
		Trees_din <= x"002f15a1";
		wait for Clk_period;
		Addr <=  "0010101100111";
		Trees_din <= x"000015a1";
		wait for Clk_period;
		Addr <=  "0010101101000";
		Trees_din <= x"13004f1c";
		wait for Clk_period;
		Addr <=  "0010101101001";
		Trees_din <= x"d4ff8710";
		wait for Clk_period;
		Addr <=  "0010101101010";
		Trees_din <= x"ebff9708";
		wait for Clk_period;
		Addr <=  "0010101101011";
		Trees_din <= x"96ffb004";
		wait for Clk_period;
		Addr <=  "0010101101100";
		Trees_din <= x"ffa51605";
		wait for Clk_period;
		Addr <=  "0010101101101";
		Trees_din <= x"00061605";
		wait for Clk_period;
		Addr <=  "0010101101110";
		Trees_din <= x"eeffcb04";
		wait for Clk_period;
		Addr <=  "0010101101111";
		Trees_din <= x"fff51605";
		wait for Clk_period;
		Addr <=  "0010101110000";
		Trees_din <= x"00561605";
		wait for Clk_period;
		Addr <=  "0010101110001";
		Trees_din <= x"93ffe108";
		wait for Clk_period;
		Addr <=  "0010101110010";
		Trees_din <= x"c8ffd304";
		wait for Clk_period;
		Addr <=  "0010101110011";
		Trees_din <= x"000f1605";
		wait for Clk_period;
		Addr <=  "0010101110100";
		Trees_din <= x"006b1605";
		wait for Clk_period;
		Addr <=  "0010101110101";
		Trees_din <= x"fffd1605";
		wait for Clk_period;
		Addr <=  "0010101110110";
		Trees_din <= x"34ffd310";
		wait for Clk_period;
		Addr <=  "0010101110111";
		Trees_din <= x"0eff5c08";
		wait for Clk_period;
		Addr <=  "0010101111000";
		Trees_din <= x"86ff8d04";
		wait for Clk_period;
		Addr <=  "0010101111001";
		Trees_din <= x"ffa61605";
		wait for Clk_period;
		Addr <=  "0010101111010";
		Trees_din <= x"00151605";
		wait for Clk_period;
		Addr <=  "0010101111011";
		Trees_din <= x"22007504";
		wait for Clk_period;
		Addr <=  "0010101111100";
		Trees_din <= x"fff91605";
		wait for Clk_period;
		Addr <=  "0010101111101";
		Trees_din <= x"005c1605";
		wait for Clk_period;
		Addr <=  "0010101111110";
		Trees_din <= x"0cffe904";
		wait for Clk_period;
		Addr <=  "0010101111111";
		Trees_din <= x"ff821605";
		wait for Clk_period;
		Addr <=  "0010110000000";
		Trees_din <= x"00011605";
		wait for Clk_period;
		Addr <=  "0010110000001";
		Trees_din <= x"70ff100c";
		wait for Clk_period;
		Addr <=  "0010110000010";
		Trees_din <= x"84008408";
		wait for Clk_period;
		Addr <=  "0010110000011";
		Trees_din <= x"04ffd704";
		wait for Clk_period;
		Addr <=  "0010110000100";
		Trees_din <= x"fff81659";
		wait for Clk_period;
		Addr <=  "0010110000101";
		Trees_din <= x"ff811659";
		wait for Clk_period;
		Addr <=  "0010110000110";
		Trees_din <= x"00221659";
		wait for Clk_period;
		Addr <=  "0010110000111";
		Trees_din <= x"85fff510";
		wait for Clk_period;
		Addr <=  "0010110001000";
		Trees_din <= x"92ffb008";
		wait for Clk_period;
		Addr <=  "0010110001001";
		Trees_din <= x"76003104";
		wait for Clk_period;
		Addr <=  "0010110001010";
		Trees_din <= x"ff9d1659";
		wait for Clk_period;
		Addr <=  "0010110001011";
		Trees_din <= x"00031659";
		wait for Clk_period;
		Addr <=  "0010110001100";
		Trees_din <= x"d2ff1604";
		wait for Clk_period;
		Addr <=  "0010110001101";
		Trees_din <= x"004b1659";
		wait for Clk_period;
		Addr <=  "0010110001110";
		Trees_din <= x"ffd41659";
		wait for Clk_period;
		Addr <=  "0010110001111";
		Trees_din <= x"0b00ad0c";
		wait for Clk_period;
		Addr <=  "0010110010000";
		Trees_din <= x"d9ffaf04";
		wait for Clk_period;
		Addr <=  "0010110010001";
		Trees_din <= x"fff61659";
		wait for Clk_period;
		Addr <=  "0010110010010";
		Trees_din <= x"34ffdd04";
		wait for Clk_period;
		Addr <=  "0010110010011";
		Trees_din <= x"00761659";
		wait for Clk_period;
		Addr <=  "0010110010100";
		Trees_din <= x"00221659";
		wait for Clk_period;
		Addr <=  "0010110010101";
		Trees_din <= x"ffdd1659";
		wait for Clk_period;
		Addr <=  "0010110010110";
		Trees_din <= x"14ff4a08";
		wait for Clk_period;
		Addr <=  "0010110010111";
		Trees_din <= x"00ffbe04";
		wait for Clk_period;
		Addr <=  "0010110011000";
		Trees_din <= x"ff8216b5";
		wait for Clk_period;
		Addr <=  "0010110011001";
		Trees_din <= x"000816b5";
		wait for Clk_period;
		Addr <=  "0010110011010";
		Trees_din <= x"96ffca18";
		wait for Clk_period;
		Addr <=  "0010110011011";
		Trees_din <= x"b8ffb508";
		wait for Clk_period;
		Addr <=  "0010110011100";
		Trees_din <= x"83ff1104";
		wait for Clk_period;
		Addr <=  "0010110011101";
		Trees_din <= x"fff716b5";
		wait for Clk_period;
		Addr <=  "0010110011110";
		Trees_din <= x"ffa016b5";
		wait for Clk_period;
		Addr <=  "0010110011111";
		Trees_din <= x"baff7c08";
		wait for Clk_period;
		Addr <=  "0010110100000";
		Trees_din <= x"e5ff0504";
		wait for Clk_period;
		Addr <=  "0010110100001";
		Trees_din <= x"001116b5";
		wait for Clk_period;
		Addr <=  "0010110100010";
		Trees_din <= x"005616b5";
		wait for Clk_period;
		Addr <=  "0010110100011";
		Trees_din <= x"24ff8704";
		wait for Clk_period;
		Addr <=  "0010110100100";
		Trees_din <= x"001316b5";
		wait for Clk_period;
		Addr <=  "0010110100101";
		Trees_din <= x"ffbc16b5";
		wait for Clk_period;
		Addr <=  "0010110100110";
		Trees_din <= x"83ff710c";
		wait for Clk_period;
		Addr <=  "0010110100111";
		Trees_din <= x"f7ff6d08";
		wait for Clk_period;
		Addr <=  "0010110101000";
		Trees_din <= x"e2ff5d04";
		wait for Clk_period;
		Addr <=  "0010110101001";
		Trees_din <= x"007316b5";
		wait for Clk_period;
		Addr <=  "0010110101010";
		Trees_din <= x"002216b5";
		wait for Clk_period;
		Addr <=  "0010110101011";
		Trees_din <= x"ffea16b5";
		wait for Clk_period;
		Addr <=  "0010110101100";
		Trees_din <= x"ffe216b5";
		wait for Clk_period;
		Addr <=  "0010110101101";
		Trees_din <= x"0eff000c";
		wait for Clk_period;
		Addr <=  "0010110101110";
		Trees_din <= x"e9ff7b04";
		wait for Clk_period;
		Addr <=  "0010110101111";
		Trees_din <= x"ff8b1711";
		wait for Clk_period;
		Addr <=  "0010110110000";
		Trees_din <= x"c1fee704";
		wait for Clk_period;
		Addr <=  "0010110110001";
		Trees_din <= x"ffcb1711";
		wait for Clk_period;
		Addr <=  "0010110110010";
		Trees_din <= x"002b1711";
		wait for Clk_period;
		Addr <=  "0010110110011";
		Trees_din <= x"b0ff6f08";
		wait for Clk_period;
		Addr <=  "0010110110100";
		Trees_din <= x"9dff5c04";
		wait for Clk_period;
		Addr <=  "0010110110101";
		Trees_din <= x"000d1711";
		wait for Clk_period;
		Addr <=  "0010110110110";
		Trees_din <= x"ffaa1711";
		wait for Clk_period;
		Addr <=  "0010110110111";
		Trees_din <= x"ba000118";
		wait for Clk_period;
		Addr <=  "0010110111000";
		Trees_din <= x"83ff3e0c";
		wait for Clk_period;
		Addr <=  "0010110111001";
		Trees_din <= x"e2ff3504";
		wait for Clk_period;
		Addr <=  "0010110111010";
		Trees_din <= x"006e1711";
		wait for Clk_period;
		Addr <=  "0010110111011";
		Trees_din <= x"48002404";
		wait for Clk_period;
		Addr <=  "0010110111100";
		Trees_din <= x"003d1711";
		wait for Clk_period;
		Addr <=  "0010110111101";
		Trees_din <= x"ffde1711";
		wait for Clk_period;
		Addr <=  "0010110111110";
		Trees_din <= x"b8ffba04";
		wait for Clk_period;
		Addr <=  "0010110111111";
		Trees_din <= x"ffbc1711";
		wait for Clk_period;
		Addr <=  "0010111000000";
		Trees_din <= x"b6ff8b04";
		wait for Clk_period;
		Addr <=  "0010111000001";
		Trees_din <= x"fff81711";
		wait for Clk_period;
		Addr <=  "0010111000010";
		Trees_din <= x"004e1711";
		wait for Clk_period;
		Addr <=  "0010111000011";
		Trees_din <= x"ffcd1711";
		wait for Clk_period;
		Addr <=  "0010111000100";
		Trees_din <= x"13004f18";
		wait for Clk_period;
		Addr <=  "0010111000101";
		Trees_din <= x"6bfeb808";
		wait for Clk_period;
		Addr <=  "0010111000110";
		Trees_din <= x"3bff1804";
		wait for Clk_period;
		Addr <=  "0010111000111";
		Trees_din <= x"00221765";
		wait for Clk_period;
		Addr <=  "0010111001000";
		Trees_din <= x"ffb51765";
		wait for Clk_period;
		Addr <=  "0010111001001";
		Trees_din <= x"96ffca0c";
		wait for Clk_period;
		Addr <=  "0010111001010";
		Trees_din <= x"e9ff8604";
		wait for Clk_period;
		Addr <=  "0010111001011";
		Trees_din <= x"ffcc1765";
		wait for Clk_period;
		Addr <=  "0010111001100";
		Trees_din <= x"a0ff3904";
		wait for Clk_period;
		Addr <=  "0010111001101";
		Trees_din <= x"00451765";
		wait for Clk_period;
		Addr <=  "0010111001110";
		Trees_din <= x"000c1765";
		wait for Clk_period;
		Addr <=  "0010111001111";
		Trees_din <= x"00591765";
		wait for Clk_period;
		Addr <=  "0010111010000";
		Trees_din <= x"34ffd30c";
		wait for Clk_period;
		Addr <=  "0010111010001";
		Trees_din <= x"57ff2d08";
		wait for Clk_period;
		Addr <=  "0010111010010";
		Trees_din <= x"0eff5c04";
		wait for Clk_period;
		Addr <=  "0010111010011";
		Trees_din <= x"fff41765";
		wait for Clk_period;
		Addr <=  "0010111010100";
		Trees_din <= x"00481765";
		wait for Clk_period;
		Addr <=  "0010111010101";
		Trees_din <= x"ffc91765";
		wait for Clk_period;
		Addr <=  "0010111010110";
		Trees_din <= x"14ffa504";
		wait for Clk_period;
		Addr <=  "0010111010111";
		Trees_din <= x"ff861765";
		wait for Clk_period;
		Addr <=  "0010111011000";
		Trees_din <= x"ffed1765";
		wait for Clk_period;
		Addr <=  "0010111011001";
		Trees_din <= x"70ff100c";
		wait for Clk_period;
		Addr <=  "0010111011010";
		Trees_din <= x"d2ff4b08";
		wait for Clk_period;
		Addr <=  "0010111011011";
		Trees_din <= x"32ff8b04";
		wait for Clk_period;
		Addr <=  "0010111011100";
		Trees_din <= x"ff8c17b9";
		wait for Clk_period;
		Addr <=  "0010111011101";
		Trees_din <= x"ffde17b9";
		wait for Clk_period;
		Addr <=  "0010111011110";
		Trees_din <= x"000d17b9";
		wait for Clk_period;
		Addr <=  "0010111011111";
		Trees_din <= x"85fff510";
		wait for Clk_period;
		Addr <=  "0010111100000";
		Trees_din <= x"92ffb008";
		wait for Clk_period;
		Addr <=  "0010111100001";
		Trees_din <= x"a3ff4804";
		wait for Clk_period;
		Addr <=  "0010111100010";
		Trees_din <= x"000017b9";
		wait for Clk_period;
		Addr <=  "0010111100011";
		Trees_din <= x"ffa317b9";
		wait for Clk_period;
		Addr <=  "0010111100100";
		Trees_din <= x"d2ff1604";
		wait for Clk_period;
		Addr <=  "0010111100101";
		Trees_din <= x"004017b9";
		wait for Clk_period;
		Addr <=  "0010111100110";
		Trees_din <= x"ffda17b9";
		wait for Clk_period;
		Addr <=  "0010111100111";
		Trees_din <= x"03ff6308";
		wait for Clk_period;
		Addr <=  "0010111101000";
		Trees_din <= x"d9ffa804";
		wait for Clk_period;
		Addr <=  "0010111101001";
		Trees_din <= x"000417b9";
		wait for Clk_period;
		Addr <=  "0010111101010";
		Trees_din <= x"006317b9";
		wait for Clk_period;
		Addr <=  "0010111101011";
		Trees_din <= x"22000504";
		wait for Clk_period;
		Addr <=  "0010111101100";
		Trees_din <= x"002917b9";
		wait for Clk_period;
		Addr <=  "0010111101101";
		Trees_din <= x"ffd317b9";
		wait for Clk_period;
		Addr <=  "0010111101110";
		Trees_din <= x"0cfeff0c";
		wait for Clk_period;
		Addr <=  "0010111101111";
		Trees_din <= x"8dfefd04";
		wait for Clk_period;
		Addr <=  "0010111110000";
		Trees_din <= x"ff8e17fd";
		wait for Clk_period;
		Addr <=  "0010111110001";
		Trees_din <= x"17001104";
		wait for Clk_period;
		Addr <=  "0010111110010";
		Trees_din <= x"ffb317fd";
		wait for Clk_period;
		Addr <=  "0010111110011";
		Trees_din <= x"003617fd";
		wait for Clk_period;
		Addr <=  "0010111110100";
		Trees_din <= x"c1feb304";
		wait for Clk_period;
		Addr <=  "0010111110101";
		Trees_din <= x"ffcc17fd";
		wait for Clk_period;
		Addr <=  "0010111110110";
		Trees_din <= x"83ff7110";
		wait for Clk_period;
		Addr <=  "0010111110111";
		Trees_din <= x"25ffdd04";
		wait for Clk_period;
		Addr <=  "0010111111000";
		Trees_din <= x"fff017fd";
		wait for Clk_period;
		Addr <=  "0010111111001";
		Trees_din <= x"e9ff2704";
		wait for Clk_period;
		Addr <=  "0010111111010";
		Trees_din <= x"000517fd";
		wait for Clk_period;
		Addr <=  "0010111111011";
		Trees_din <= x"e2ff5804";
		wait for Clk_period;
		Addr <=  "0010111111100";
		Trees_din <= x"006c17fd";
		wait for Clk_period;
		Addr <=  "0010111111101";
		Trees_din <= x"001317fd";
		wait for Clk_period;
		Addr <=  "0010111111110";
		Trees_din <= x"ffdf17fd";
		wait for Clk_period;
		Addr <=  "0010111111111";
		Trees_din <= x"0eff000c";
		wait for Clk_period;
		Addr <=  "0011000000000";
		Trees_din <= x"0cffc208";
		wait for Clk_period;
		Addr <=  "0011000000001";
		Trees_din <= x"fcff8904";
		wait for Clk_period;
		Addr <=  "0011000000010";
		Trees_din <= x"ff8f1851";
		wait for Clk_period;
		Addr <=  "0011000000011";
		Trees_din <= x"ffeb1851";
		wait for Clk_period;
		Addr <=  "0011000000100";
		Trees_din <= x"00161851";
		wait for Clk_period;
		Addr <=  "0011000000101";
		Trees_din <= x"75009e18";
		wait for Clk_period;
		Addr <=  "0011000000110";
		Trees_din <= x"dfffb510";
		wait for Clk_period;
		Addr <=  "0011000000111";
		Trees_din <= x"81ff7408";
		wait for Clk_period;
		Addr <=  "0011000001000";
		Trees_din <= x"da003104";
		wait for Clk_period;
		Addr <=  "0011000001001";
		Trees_din <= x"ffe71851";
		wait for Clk_period;
		Addr <=  "0011000001010";
		Trees_din <= x"003f1851";
		wait for Clk_period;
		Addr <=  "0011000001011";
		Trees_din <= x"9dff4f04";
		wait for Clk_period;
		Addr <=  "0011000001100";
		Trees_din <= x"000f1851";
		wait for Clk_period;
		Addr <=  "0011000001101";
		Trees_din <= x"ffab1851";
		wait for Clk_period;
		Addr <=  "0011000001110";
		Trees_din <= x"b6ff9504";
		wait for Clk_period;
		Addr <=  "0011000001111";
		Trees_din <= x"00021851";
		wait for Clk_period;
		Addr <=  "0011000010000";
		Trees_din <= x"00451851";
		wait for Clk_period;
		Addr <=  "0011000010001";
		Trees_din <= x"baff9f04";
		wait for Clk_period;
		Addr <=  "0011000010010";
		Trees_din <= x"00561851";
		wait for Clk_period;
		Addr <=  "0011000010011";
		Trees_din <= x"00141851";
		wait for Clk_period;
		Addr <=  "0011000010100";
		Trees_din <= x"1300d518";
		wait for Clk_period;
		Addr <=  "0011000010101";
		Trees_din <= x"b0ff6104";
		wait for Clk_period;
		Addr <=  "0011000010110";
		Trees_din <= x"ffbc1885";
		wait for Clk_period;
		Addr <=  "0011000010111";
		Trees_din <= x"b8ff5a04";
		wait for Clk_period;
		Addr <=  "0011000011000";
		Trees_din <= x"ffd31885";
		wait for Clk_period;
		Addr <=  "0011000011001";
		Trees_din <= x"57ff820c";
		wait for Clk_period;
		Addr <=  "0011000011010";
		Trees_din <= x"9fff2604";
		wait for Clk_period;
		Addr <=  "0011000011011";
		Trees_din <= x"fff11885";
		wait for Clk_period;
		Addr <=  "0011000011100";
		Trees_din <= x"c1feb204";
		wait for Clk_period;
		Addr <=  "0011000011101";
		Trees_din <= x"fff71885";
		wait for Clk_period;
		Addr <=  "0011000011110";
		Trees_din <= x"00551885";
		wait for Clk_period;
		Addr <=  "0011000011111";
		Trees_din <= x"ffe21885";
		wait for Clk_period;
		Addr <=  "0011000100000";
		Trees_din <= x"ffa81885";
		wait for Clk_period;
		Addr <=  "0011000100001";
		Trees_din <= x"70ff240c";
		wait for Clk_period;
		Addr <=  "0011000100010";
		Trees_din <= x"ebff6008";
		wait for Clk_period;
		Addr <=  "0011000100011";
		Trees_din <= x"c7ff6b04";
		wait for Clk_period;
		Addr <=  "0011000100100";
		Trees_din <= x"ff9618c9";
		wait for Clk_period;
		Addr <=  "0011000100101";
		Trees_din <= x"ffe518c9";
		wait for Clk_period;
		Addr <=  "0011000100110";
		Trees_din <= x"000d18c9";
		wait for Clk_period;
		Addr <=  "0011000100111";
		Trees_din <= x"85fff50c";
		wait for Clk_period;
		Addr <=  "0011000101000";
		Trees_din <= x"baff6704";
		wait for Clk_period;
		Addr <=  "0011000101001";
		Trees_din <= x"002a18c9";
		wait for Clk_period;
		Addr <=  "0011000101010";
		Trees_din <= x"51000204";
		wait for Clk_period;
		Addr <=  "0011000101011";
		Trees_din <= x"ffb218c9";
		wait for Clk_period;
		Addr <=  "0011000101100";
		Trees_din <= x"001218c9";
		wait for Clk_period;
		Addr <=  "0011000101101";
		Trees_din <= x"03ff8308";
		wait for Clk_period;
		Addr <=  "0011000101110";
		Trees_din <= x"4fff9c04";
		wait for Clk_period;
		Addr <=  "0011000101111";
		Trees_din <= x"000f18c9";
		wait for Clk_period;
		Addr <=  "0011000110000";
		Trees_din <= x"005a18c9";
		wait for Clk_period;
		Addr <=  "0011000110001";
		Trees_din <= x"fff618c9";
		wait for Clk_period;
		Addr <=  "0011000110010";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  4
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"51010650";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"89015538";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"8e00f020";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"8a004310";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"5100c908";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"c2005e04";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"ff6a00fd";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"000b00fd";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"fb003604";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"ffc900fd";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"01d200fd";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"90006708";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"9ffe9b04";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"019a00fd";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"ff9600fd";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"e8ffc504";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"023d00fd";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"ff7c00fd";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"64ff050c";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"5a008c08";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"0ffedb04";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"032f00fd";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"00ca00fd";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"000000fd";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"69ff8c04";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"ff6500fd";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"33ff5304";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"ff9c00fd";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"01ef00fd";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"1f00a010";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"d4fefb08";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"00ffaf04";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"ff9000fd";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"003700fd";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"12ffb804";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"008900fd";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"03d400fd";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"90ffda04";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"ff6800fd";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"01b000fd";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"90fffb1c";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"faff920c";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"78fefd08";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"18ff9204";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"015c00fd";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"ff9000fd";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"ff5e00fd";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"11ff7804";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"ff7c00fd";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"7d001b04";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"033300fd";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"04009304";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"00ca00fd";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"ff9600fd";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"a3ff2a04";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"ff9600fd";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"f3fe3d04";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"ffa400fd";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"8dfdf404";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"003700fd";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"56ff8804";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"042f00fd";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"00ca00fd";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"5100d15c";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"8900be28";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"8e01231c";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"0b014910";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"a3ffa908";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"bffe2004";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"00050239";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"ff660239";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"8a007004";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"ff8e0239";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"007c0239";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"deff6008";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"17ff9604";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"00260239";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"023f0239";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"ff7b0239";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"aaff5504";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"ff7f0239";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"a7ffa604";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"00020239";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"02190239";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"8e001d1c";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"d5ffad0c";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"23000104";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"ff850239";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"92fec704";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"00250239";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"02850239";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"cfffea08";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"c2000604";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"ff740239";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"01bc0239";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"7ffdb204";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"00ac0239";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"ff630239";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"00ff8608";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"05002304";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"014c0239";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"ff670239";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"83ff5008";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"06fed304";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"fff20239";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"02250239";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"14ff0304";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"ff860239";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"003a0239";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"8dfe8c1c";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"a9fee310";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"baff9c08";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"70fe7704";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"002e0239";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"02240239";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"67ff1004";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"00390239";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"ff8c0239";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"ddfe2204";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"01120239";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"bf001504";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"ff5a0239";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"006f0239";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"2fffe114";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"5bff2204";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"ff6f0239";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"22004c08";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"7d001004";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"01cb0239";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"002f0239";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"5bff6204";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"003c0239";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"ff870239";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"15ffee10";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"8c00b608";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"bcffa204";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"02260239";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"00200239";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"0cfde904";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"01170239";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"ff910239";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"ff9c0239";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"8a004370";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"5100c93c";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"8900f420";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"8e00f010";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"7fffe608";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"43005504";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"ff6f03a5";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"001203a5";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"39ff9a04";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"001003a5";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"ff7403a5";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"7fffa808";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"feff3b04";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"00ba03a5";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"ff6b03a5";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"58feda04";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"019703a5";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"002403a5";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"b6ff5a10";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"6aff9808";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"6fff4104";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"01bd03a5";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"ffa603a5";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"6d004a04";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"ff8503a5";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"003003a5";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"e5ff3408";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"b3ff7904";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"ff6303a5";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"002803a5";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"00b203a5";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"efff5714";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"7bff7910";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"96ff0308";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"05006404";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"002403a5";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"ffa603a5";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"c0ff7304";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"01df03a5";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"000b03a5";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"ff9403a5";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"69fe6910";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"70feca08";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"dfff2a04";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"006703a5";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"019303a5";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"d9ffd204";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"003003a5";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"ff9f03a5";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"b0ff9308";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"89009e04";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"ff5c03a5";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"003103a5";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"9eff7f04";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"012e03a5";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"ff8a03a5";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"e4fe2c24";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"4bff4218";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"0dff380c";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"64ff5708";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"b6feef04";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"009703a5";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"01bd03a5";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"ff9e03a5";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"8a00b604";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"ff7403a5";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"43ff4f04";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"001e03a5";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"014703a5";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"64fe9d08";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"32fecc04";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"014503a5";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"ffa203a5";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"ff6c03a5";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"30008b18";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"16fdde08";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"32fe9504";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"019e03a5";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"ff9d03a5";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"1effe108";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"b8fe6304";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"003d03a5";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"ff6a03a5";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"69ff0f04";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"014903a5";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"ff7403a5";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"efffb408";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"b2fff004";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"01eb03a5";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"002c03a5";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"ffa203a5";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"8a00435c";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"dc00b734";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"8900f41c";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"b7febc0c";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"a1fedf04";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"ff7204e9";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"1afeb604";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"01bd04e9";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"ffde04e9";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"7fffe608";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"43005504";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"ff7404e9";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"001804e9";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"c5ff3104";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"002704e9";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"ff7004e9";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"6aff9810";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"c2000008";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"0a00e004";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"ff9704e9";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"00c104e9";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"efff8904";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"01a604e9";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"002004e9";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"8e00d604";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"ff6804e9";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"009504e9";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"faff6e0c";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"28ffc004";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"ff6304e9";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"8e003b04";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"ffab04e9";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"013e04e9";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"30ffd40c";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"c5ff0e08";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"67fe8104";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"010d04e9";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"000004e9";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"ff7004e9";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"fdff2908";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"ab00c404";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"ff8f04e9";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"003204e9";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"c6ff1b04";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"01f104e9";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"000b04e9";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"e4fe2c1c";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"98fe3704";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"ff7c04e9";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"2200280c";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"a7010108";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"1f00fc04";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"012d04e9";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"ff9904e9";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"ff9204e9";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"9bff0d08";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"72ffe304";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"011b04e9";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"001704e9";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"ff7704e9";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"30008b20";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"e9fe8010";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"a3ffa108";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"85ff3004";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"008e04e9";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"ff6c04e9";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"f9fea804";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"ff9404e9";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"012d04e9";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"8e009508";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"88015404";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"ff6a04e9";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"008d04e9";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"4aff5e04";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"00cb04e9";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"002304e9";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"efffb408";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"7bff0504";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"016f04e9";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"002304e9";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"ffa804e9";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"8a004370";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"2fffec40";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"00ffe120";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"1cfec610";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"0fff2f08";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"7affa704";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"ffdd064d";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"020b064d";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"62ffae04";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"ff8b064d";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"014a064d";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"8e00d608";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"88014004";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"ff74064d";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"0024064d";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"50ff0a04";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"0108064d";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"ff97064d";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"6fff4710";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"62ff6f08";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"88003f04";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"ffb7064d";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"00e4064d";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"66ffd304";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"0040064d";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"02b9064d";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"5100ba08";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"d9002804";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"ff67064d";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"0047064d";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"67fedf04";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"00fe064d";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"0007064d";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"c5ff1714";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"1eff9e04";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"ff82064d";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"70ff2608";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"8dfee804";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"ffe0064d";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"0132064d";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"06ff4604";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"0073064d";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"0353064d";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"73003d10";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"40ff9a08";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"04005704";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"ffa6064d";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"0160064d";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"a7ff5b04";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"0001064d";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"ff66064d";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"17ffdf04";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"ff7d064d";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"0efe9e04";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"ff95064d";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"0155064d";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"e4fe161c";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"4bff4210";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"00ff1004";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"ff97064d";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"de00b008";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"64ff5704";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"010f064d";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"fff9064d";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"ff96064d";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"68fec708";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"08006b04";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"00c9064d";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"fff9064d";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"ff75064d";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"bfff0d14";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"0800bf0c";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"82ff6808";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"4f005104";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"0115064d";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"ffd6064d";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"ff92064d";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"6aff3904";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"0028064d";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"ff76064d";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"84015b10";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"74004108";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"28ffcf04";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"ff6d064d";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"006c064d";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"eaff9604";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"ff7e064d";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"00f2064d";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"00d0064d";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"0a00443c";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"43fe720c";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"87ff6304";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"ff9807a1";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"01fe9304";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"002007a1";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"01e507a1";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"ccff0618";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"a9ff1e0c";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"7c001b08";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"d7007904";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"ff9307a1";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"009b07a1";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"01fe07a1";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"5efeb004";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"012607a1";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"0a003704";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"ff6607a1";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"009007a1";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"2e00a810";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"40ff8008";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"f202ec04";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"ff8207a1";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"016407a1";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"8900f404";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"ff7207a1";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"001407a1";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"8aff7e04";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"ffaf07a1";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"014e07a1";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"67ff7240";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"c3ffb820";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"8dfe9610";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"7d003808";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"b2004904";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"ff6c07a1";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"008507a1";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"d000af04";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"ffcd07a1";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"010307a1";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"14ff6d08";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"b8ff2704";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"007907a1";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"015807a1";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"ccfee104";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"008807a1";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"ff7a07a1";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"90ffe610";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"84009008";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"3cfe7e04";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"00ca07a1";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"ffa307a1";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"51005004";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"ffc107a1";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"00e707a1";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"89008a08";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"fb006004";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"ffc407a1";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"011a07a1";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"4aff7104";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"012607a1";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"fffb07a1";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"b5fe6014";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"a7ff9804";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"ff7a07a1";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"30ffc108";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"2dfe9e04";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"fff607a1";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"ff9807a1";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"40003c04";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"013807a1";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"ff9d07a1";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"42fffe0c";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"43007308";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"46fe3d04";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"fff507a1";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"ff6207a1";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"008a07a1";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"adffcd08";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"51ff4f04";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"003807a1";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"ff6e07a1";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"86ff4a04";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"ffe507a1";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"016707a1";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"0a00464c";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"ccff2c28";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"9c00021c";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"f0febf0c";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"fdffa204";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"ffae08fd";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"2cff8504";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"01ef08fd";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"007908fd";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"19fed408";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"fdff6e04";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"ffa508fd";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"010908fd";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"10010504";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"ff6508fd";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"003c08fd";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"f2021204";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"ffa108fd";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"74ffe104";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"000d08fd";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"018f08fd";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"43fe7208";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"aaff8904";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"ffa008fd";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"012008fd";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"00ffde0c";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"b3fff808";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"40ff6304";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"009108fd";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"ff7208fd";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"00b608fd";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"3d000808";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"5dff4004";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"004308fd";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"ff6f08fd";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"f6fee304";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"ff9508fd";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"010c08fd";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"67ff7234";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"11ff8f14";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"d3fe1e04";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"016308fd";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"89002f08";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"74003c04";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"ff7808fd";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"001e08fd";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"7dff3e04";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"016708fd";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"fff608fd";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"39ffb210";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"73ffd008";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"b5ff0b04";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"006108fd";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"ff7408fd";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"34003a04";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"00e308fd";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"ffb808fd";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"c3ffdf08";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"a1ff0004";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"ffab08fd";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"008908fd";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"9afe7504";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"001c08fd";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"ff6908fd";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"b5fe6014";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"a7ff9804";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"ff8008fd";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"63ff6e08";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"b9fea504";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"ffea08fd";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"012e08fd";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"1b00fc04";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"ff8808fd";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"007c08fd";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"42fffe0c";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"43007308";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"81fef104";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"000408fd";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"ff6508fd";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"007908fd";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"ceff8b08";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"f2020404";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"012408fd";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"ffef08fd";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"dffec904";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"002608fd";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"ff7308fd";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"0a00464c";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"9cff9420";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"2e00a818";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"43fe8d0c";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"58fe7e08";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"8e001104";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"00120a61";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"00f90a61";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"ff930a61";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"50008908";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"88ff1804";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"002b0a61";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"ff6c0a61";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"00650a61";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"d6006b04";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"00c60a61";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"00230a61";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"5fffc720";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"0fff2910";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"aaffed08";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"ccff2404";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"00b90a61";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"ff730a61";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"c8000304";
		wait for Clk_period;
		Addr <=  "0001001010111";
		Trees_din <= x"00350a61";
		wait for Clk_period;
		Addr <=  "0001001011000";
		Trees_din <= x"02050a61";
		wait for Clk_period;
		Addr <=  "0001001011001";
		Trees_din <= x"40ff8b08";
		wait for Clk_period;
		Addr <=  "0001001011010";
		Trees_din <= x"a3ffa404";
		wait for Clk_period;
		Addr <=  "0001001011011";
		Trees_din <= x"ff950a61";
		wait for Clk_period;
		Addr <=  "0001001011100";
		Trees_din <= x"01520a61";
		wait for Clk_period;
		Addr <=  "0001001011101";
		Trees_din <= x"c5fec604";
		wait for Clk_period;
		Addr <=  "0001001011110";
		Trees_din <= x"00a50a61";
		wait for Clk_period;
		Addr <=  "0001001011111";
		Trees_din <= x"ff7c0a61";
		wait for Clk_period;
		Addr <=  "0001001100000";
		Trees_din <= x"12ff7c04";
		wait for Clk_period;
		Addr <=  "0001001100001";
		Trees_din <= x"ff880a61";
		wait for Clk_period;
		Addr <=  "0001001100010";
		Trees_din <= x"4cff3c04";
		wait for Clk_period;
		Addr <=  "0001001100011";
		Trees_din <= x"023e0a61";
		wait for Clk_period;
		Addr <=  "0001001100100";
		Trees_din <= x"00590a61";
		wait for Clk_period;
		Addr <=  "0001001100101";
		Trees_din <= x"0fff2f34";
		wait for Clk_period;
		Addr <=  "0001001100110";
		Trees_din <= x"aaff7818";
		wait for Clk_period;
		Addr <=  "0001001100111";
		Trees_din <= x"88001c08";
		wait for Clk_period;
		Addr <=  "0001001101000";
		Trees_din <= x"58fe5004";
		wait for Clk_period;
		Addr <=  "0001001101001";
		Trees_din <= x"00380a61";
		wait for Clk_period;
		Addr <=  "0001001101010";
		Trees_din <= x"ff6a0a61";
		wait for Clk_period;
		Addr <=  "0001001101011";
		Trees_din <= x"cafe7508";
		wait for Clk_period;
		Addr <=  "0001001101100";
		Trees_din <= x"0a008404";
		wait for Clk_period;
		Addr <=  "0001001101101";
		Trees_din <= x"ffbf0a61";
		wait for Clk_period;
		Addr <=  "0001001101110";
		Trees_din <= x"00b90a61";
		wait for Clk_period;
		Addr <=  "0001001101111";
		Trees_din <= x"6aff1f04";
		wait for Clk_period;
		Addr <=  "0001001110000";
		Trees_din <= x"00720a61";
		wait for Clk_period;
		Addr <=  "0001001110001";
		Trees_din <= x"ff850a61";
		wait for Clk_period;
		Addr <=  "0001001110010";
		Trees_din <= x"c3ffea10";
		wait for Clk_period;
		Addr <=  "0001001110011";
		Trees_din <= x"17ff9208";
		wait for Clk_period;
		Addr <=  "0001001110100";
		Trees_din <= x"84007004";
		wait for Clk_period;
		Addr <=  "0001001110101";
		Trees_din <= x"ff910a61";
		wait for Clk_period;
		Addr <=  "0001001110110";
		Trees_din <= x"00540a61";
		wait for Clk_period;
		Addr <=  "0001001110111";
		Trees_din <= x"5a00c804";
		wait for Clk_period;
		Addr <=  "0001001111000";
		Trees_din <= x"01150a61";
		wait for Clk_period;
		Addr <=  "0001001111001";
		Trees_din <= x"00240a61";
		wait for Clk_period;
		Addr <=  "0001001111010";
		Trees_din <= x"69ff3608";
		wait for Clk_period;
		Addr <=  "0001001111011";
		Trees_din <= x"79ff4604";
		wait for Clk_period;
		Addr <=  "0001001111100";
		Trees_din <= x"00080a61";
		wait for Clk_period;
		Addr <=  "0001001111101";
		Trees_din <= x"00d30a61";
		wait for Clk_period;
		Addr <=  "0001001111110";
		Trees_din <= x"ff7a0a61";
		wait for Clk_period;
		Addr <=  "0001001111111";
		Trees_din <= x"fa000b20";
		wait for Clk_period;
		Addr <=  "0001010000000";
		Trees_din <= x"d000d810";
		wait for Clk_period;
		Addr <=  "0001010000001";
		Trees_din <= x"51010608";
		wait for Clk_period;
		Addr <=  "0001010000010";
		Trees_din <= x"bfff0904";
		wait for Clk_period;
		Addr <=  "0001010000011";
		Trees_din <= x"ffe50a61";
		wait for Clk_period;
		Addr <=  "0001010000100";
		Trees_din <= x"ff770a61";
		wait for Clk_period;
		Addr <=  "0001010000101";
		Trees_din <= x"3bff2f04";
		wait for Clk_period;
		Addr <=  "0001010000110";
		Trees_din <= x"009e0a61";
		wait for Clk_period;
		Addr <=  "0001010000111";
		Trees_din <= x"ff950a61";
		wait for Clk_period;
		Addr <=  "0001010001000";
		Trees_din <= x"37ff7908";
		wait for Clk_period;
		Addr <=  "0001010001001";
		Trees_din <= x"1eff9904";
		wait for Clk_period;
		Addr <=  "0001010001010";
		Trees_din <= x"ffce0a61";
		wait for Clk_period;
		Addr <=  "0001010001011";
		Trees_din <= x"01020a61";
		wait for Clk_period;
		Addr <=  "0001010001100";
		Trees_din <= x"87ffd504";
		wait for Clk_period;
		Addr <=  "0001010001101";
		Trees_din <= x"ff820a61";
		wait for Clk_period;
		Addr <=  "0001010001110";
		Trees_din <= x"009e0a61";
		wait for Clk_period;
		Addr <=  "0001010001111";
		Trees_din <= x"64ff3510";
		wait for Clk_period;
		Addr <=  "0001010010000";
		Trees_din <= x"3eff5508";
		wait for Clk_period;
		Addr <=  "0001010010001";
		Trees_din <= x"0cfe7404";
		wait for Clk_period;
		Addr <=  "0001010010010";
		Trees_din <= x"00350a61";
		wait for Clk_period;
		Addr <=  "0001010010011";
		Trees_din <= x"ffae0a61";
		wait for Clk_period;
		Addr <=  "0001010010100";
		Trees_din <= x"dfff7304";
		wait for Clk_period;
		Addr <=  "0001010010101";
		Trees_din <= x"00730a61";
		wait for Clk_period;
		Addr <=  "0001010010110";
		Trees_din <= x"01dc0a61";
		wait for Clk_period;
		Addr <=  "0001010010111";
		Trees_din <= x"ff890a61";
		wait for Clk_period;
		Addr <=  "0001010011000";
		Trees_din <= x"0a004344";
		wait for Clk_period;
		Addr <=  "0001010011001";
		Trees_din <= x"9cff9424";
		wait for Clk_period;
		Addr <=  "0001010011010";
		Trees_din <= x"2e00a81c";
		wait for Clk_period;
		Addr <=  "0001010011011";
		Trees_din <= x"43feac10";
		wait for Clk_period;
		Addr <=  "0001010011100";
		Trees_din <= x"aaffcc08";
		wait for Clk_period;
		Addr <=  "0001010011101";
		Trees_din <= x"8c007c04";
		wait for Clk_period;
		Addr <=  "0001010011110";
		Trees_din <= x"ff850b85";
		wait for Clk_period;
		Addr <=  "0001010011111";
		Trees_din <= x"00160b85";
		wait for Clk_period;
		Addr <=  "0001010100000";
		Trees_din <= x"f4ff2104";
		wait for Clk_period;
		Addr <=  "0001010100001";
		Trees_din <= x"ffff0b85";
		wait for Clk_period;
		Addr <=  "0001010100010";
		Trees_din <= x"01120b85";
		wait for Clk_period;
		Addr <=  "0001010100011";
		Trees_din <= x"50008908";
		wait for Clk_period;
		Addr <=  "0001010100100";
		Trees_din <= x"69fe4b04";
		wait for Clk_period;
		Addr <=  "0001010100101";
		Trees_din <= x"001d0b85";
		wait for Clk_period;
		Addr <=  "0001010100110";
		Trees_din <= x"ff6d0b85";
		wait for Clk_period;
		Addr <=  "0001010100111";
		Trees_din <= x"005d0b85";
		wait for Clk_period;
		Addr <=  "0001010101000";
		Trees_din <= x"d7005204";
		wait for Clk_period;
		Addr <=  "0001010101001";
		Trees_din <= x"001b0b85";
		wait for Clk_period;
		Addr <=  "0001010101010";
		Trees_din <= x"00c20b85";
		wait for Clk_period;
		Addr <=  "0001010101011";
		Trees_din <= x"eeff590c";
		wait for Clk_period;
		Addr <=  "0001010101100";
		Trees_din <= x"e1ffd604";
		wait for Clk_period;
		Addr <=  "0001010101101";
		Trees_din <= x"ff9a0b85";
		wait for Clk_period;
		Addr <=  "0001010101110";
		Trees_din <= x"4cff1d04";
		wait for Clk_period;
		Addr <=  "0001010101111";
		Trees_din <= x"02400b85";
		wait for Clk_period;
		Addr <=  "0001010110000";
		Trees_din <= x"00360b85";
		wait for Clk_period;
		Addr <=  "0001010110001";
		Trees_din <= x"6a00320c";
		wait for Clk_period;
		Addr <=  "0001010110010";
		Trees_din <= x"c4fdf704";
		wait for Clk_period;
		Addr <=  "0001010110011";
		Trees_din <= x"011a0b85";
		wait for Clk_period;
		Addr <=  "0001010110100";
		Trees_din <= x"5fffd704";
		wait for Clk_period;
		Addr <=  "0001010110101";
		Trees_din <= x"ff930b85";
		wait for Clk_period;
		Addr <=  "0001010110110";
		Trees_din <= x"006d0b85";
		wait for Clk_period;
		Addr <=  "0001010110111";
		Trees_din <= x"04fff804";
		wait for Clk_period;
		Addr <=  "0001010111000";
		Trees_din <= x"01c00b85";
		wait for Clk_period;
		Addr <=  "0001010111001";
		Trees_din <= x"ffa00b85";
		wait for Clk_period;
		Addr <=  "0001010111010";
		Trees_din <= x"67ff7234";
		wait for Clk_period;
		Addr <=  "0001010111011";
		Trees_din <= x"11ff7d14";
		wait for Clk_period;
		Addr <=  "0001010111100";
		Trees_din <= x"d3fe1e04";
		wait for Clk_period;
		Addr <=  "0001010111101";
		Trees_din <= x"01240b85";
		wait for Clk_period;
		Addr <=  "0001010111110";
		Trees_din <= x"3cfe9308";
		wait for Clk_period;
		Addr <=  "0001010111111";
		Trees_din <= x"2200f804";
		wait for Clk_period;
		Addr <=  "0001011000000";
		Trees_din <= x"fffc0b85";
		wait for Clk_period;
		Addr <=  "0001011000001";
		Trees_din <= x"01a80b85";
		wait for Clk_period;
		Addr <=  "0001011000010";
		Trees_din <= x"84007f04";
		wait for Clk_period;
		Addr <=  "0001011000011";
		Trees_din <= x"ff990b85";
		wait for Clk_period;
		Addr <=  "0001011000100";
		Trees_din <= x"007b0b85";
		wait for Clk_period;
		Addr <=  "0001011000101";
		Trees_din <= x"2cff7610";
		wait for Clk_period;
		Addr <=  "0001011000110";
		Trees_din <= x"dc00a508";
		wait for Clk_period;
		Addr <=  "0001011000111";
		Trees_din <= x"9efeff04";
		wait for Clk_period;
		Addr <=  "0001011001000";
		Trees_din <= x"00330b85";
		wait for Clk_period;
		Addr <=  "0001011001001";
		Trees_din <= x"ff730b85";
		wait for Clk_period;
		Addr <=  "0001011001010";
		Trees_din <= x"19ff5704";
		wait for Clk_period;
		Addr <=  "0001011001011";
		Trees_din <= x"009c0b85";
		wait for Clk_period;
		Addr <=  "0001011001100";
		Trees_din <= x"ffa50b85";
		wait for Clk_period;
		Addr <=  "0001011001101";
		Trees_din <= x"14ff7108";
		wait for Clk_period;
		Addr <=  "0001011001110";
		Trees_din <= x"39fff104";
		wait for Clk_period;
		Addr <=  "0001011001111";
		Trees_din <= x"00a30b85";
		wait for Clk_period;
		Addr <=  "0001011010000";
		Trees_din <= x"ffef0b85";
		wait for Clk_period;
		Addr <=  "0001011010001";
		Trees_din <= x"b1fe9004";
		wait for Clk_period;
		Addr <=  "0001011010010";
		Trees_din <= x"00bf0b85";
		wait for Clk_period;
		Addr <=  "0001011010011";
		Trees_din <= x"ff8c0b85";
		wait for Clk_period;
		Addr <=  "0001011010100";
		Trees_din <= x"b5fdfd08";
		wait for Clk_period;
		Addr <=  "0001011010101";
		Trees_din <= x"69ff1904";
		wait for Clk_period;
		Addr <=  "0001011010110";
		Trees_din <= x"00dd0b85";
		wait for Clk_period;
		Addr <=  "0001011010111";
		Trees_din <= x"ffe40b85";
		wait for Clk_period;
		Addr <=  "0001011011000";
		Trees_din <= x"8dffdd10";
		wait for Clk_period;
		Addr <=  "0001011011001";
		Trees_din <= x"43005508";
		wait for Clk_period;
		Addr <=  "0001011011010";
		Trees_din <= x"53fe9704";
		wait for Clk_period;
		Addr <=  "0001011011011";
		Trees_din <= x"00a00b85";
		wait for Clk_period;
		Addr <=  "0001011011100";
		Trees_din <= x"ff830b85";
		wait for Clk_period;
		Addr <=  "0001011011101";
		Trees_din <= x"b6ff4b04";
		wait for Clk_period;
		Addr <=  "0001011011110";
		Trees_din <= x"00fc0b85";
		wait for Clk_period;
		Addr <=  "0001011011111";
		Trees_din <= x"ffa50b85";
		wait for Clk_period;
		Addr <=  "0001011100000";
		Trees_din <= x"00ab0b85";
		wait for Clk_period;
		Addr <=  "0001011100001";
		Trees_din <= x"0fff314c";
		wait for Clk_period;
		Addr <=  "0001011100010";
		Trees_din <= x"1cfee11c";
		wait for Clk_period;
		Addr <=  "0001011100011";
		Trees_din <= x"78ff5910";
		wait for Clk_period;
		Addr <=  "0001011100100";
		Trees_din <= x"de00510c";
		wait for Clk_period;
		Addr <=  "0001011100101";
		Trees_din <= x"fbff5504";
		wait for Clk_period;
		Addr <=  "0001011100110";
		Trees_din <= x"fff50cc9";
		wait for Clk_period;
		Addr <=  "0001011100111";
		Trees_din <= x"a1fed704";
		wait for Clk_period;
		Addr <=  "0001011101000";
		Trees_din <= x"00380cc9";
		wait for Clk_period;
		Addr <=  "0001011101001";
		Trees_din <= x"01670cc9";
		wait for Clk_period;
		Addr <=  "0001011101010";
		Trees_din <= x"ffe70cc9";
		wait for Clk_period;
		Addr <=  "0001011101011";
		Trees_din <= x"00ff9e04";
		wait for Clk_period;
		Addr <=  "0001011101100";
		Trees_din <= x"ff8e0cc9";
		wait for Clk_period;
		Addr <=  "0001011101101";
		Trees_din <= x"6cff4304";
		wait for Clk_period;
		Addr <=  "0001011101110";
		Trees_din <= x"ffe10cc9";
		wait for Clk_period;
		Addr <=  "0001011101111";
		Trees_din <= x"00c50cc9";
		wait for Clk_period;
		Addr <=  "0001011110000";
		Trees_din <= x"c6ff2d18";
		wait for Clk_period;
		Addr <=  "0001011110001";
		Trees_din <= x"90ff6208";
		wait for Clk_period;
		Addr <=  "0001011110010";
		Trees_din <= x"4dff9f04";
		wait for Clk_period;
		Addr <=  "0001011110011";
		Trees_din <= x"ff700cc9";
		wait for Clk_period;
		Addr <=  "0001011110100";
		Trees_din <= x"00820cc9";
		wait for Clk_period;
		Addr <=  "0001011110101";
		Trees_din <= x"67ff7a08";
		wait for Clk_period;
		Addr <=  "0001011110110";
		Trees_din <= x"a7ff3e04";
		wait for Clk_period;
		Addr <=  "0001011110111";
		Trees_din <= x"ff910cc9";
		wait for Clk_period;
		Addr <=  "0001011111000";
		Trees_din <= x"00a90cc9";
		wait for Clk_period;
		Addr <=  "0001011111001";
		Trees_din <= x"b4fe6d04";
		wait for Clk_period;
		Addr <=  "0001011111010";
		Trees_din <= x"00430cc9";
		wait for Clk_period;
		Addr <=  "0001011111011";
		Trees_din <= x"ff7b0cc9";
		wait for Clk_period;
		Addr <=  "0001011111100";
		Trees_din <= x"db00f70c";
		wait for Clk_period;
		Addr <=  "0001011111101";
		Trees_din <= x"02fde804";
		wait for Clk_period;
		Addr <=  "0001011111110";
		Trees_din <= x"00ca0cc9";
		wait for Clk_period;
		Addr <=  "0001011111111";
		Trees_din <= x"7cfefb04";
		wait for Clk_period;
		Addr <=  "0001100000000";
		Trees_din <= x"00130cc9";
		wait for Clk_period;
		Addr <=  "0001100000001";
		Trees_din <= x"ff6c0cc9";
		wait for Clk_period;
		Addr <=  "0001100000010";
		Trees_din <= x"1cff8c08";
		wait for Clk_period;
		Addr <=  "0001100000011";
		Trees_din <= x"96ff2c04";
		wait for Clk_period;
		Addr <=  "0001100000100";
		Trees_din <= x"01120cc9";
		wait for Clk_period;
		Addr <=  "0001100000101";
		Trees_din <= x"00300cc9";
		wait for Clk_period;
		Addr <=  "0001100000110";
		Trees_din <= x"ff8f0cc9";
		wait for Clk_period;
		Addr <=  "0001100000111";
		Trees_din <= x"30ffb51c";
		wait for Clk_period;
		Addr <=  "0001100001000";
		Trees_din <= x"2c006810";
		wait for Clk_period;
		Addr <=  "0001100001001";
		Trees_din <= x"5101630c";
		wait for Clk_period;
		Addr <=  "0001100001010";
		Trees_din <= x"35001608";
		wait for Clk_period;
		Addr <=  "0001100001011";
		Trees_din <= x"79fe8104";
		wait for Clk_period;
		Addr <=  "0001100001100";
		Trees_din <= x"fff60cc9";
		wait for Clk_period;
		Addr <=  "0001100001101";
		Trees_din <= x"ff620cc9";
		wait for Clk_period;
		Addr <=  "0001100001110";
		Trees_din <= x"00210cc9";
		wait for Clk_period;
		Addr <=  "0001100001111";
		Trees_din <= x"005b0cc9";
		wait for Clk_period;
		Addr <=  "0001100010000";
		Trees_din <= x"50ff1f08";
		wait for Clk_period;
		Addr <=  "0001100010001";
		Trees_din <= x"02fe4704";
		wait for Clk_period;
		Addr <=  "0001100010010";
		Trees_din <= x"01650cc9";
		wait for Clk_period;
		Addr <=  "0001100010011";
		Trees_din <= x"00500cc9";
		wait for Clk_period;
		Addr <=  "0001100010100";
		Trees_din <= x"ff900cc9";
		wait for Clk_period;
		Addr <=  "0001100010101";
		Trees_din <= x"faffc820";
		wait for Clk_period;
		Addr <=  "0001100010110";
		Trees_din <= x"1afecf10";
		wait for Clk_period;
		Addr <=  "0001100010111";
		Trees_din <= x"ebfee308";
		wait for Clk_period;
		Addr <=  "0001100011000";
		Trees_din <= x"00ffc304";
		wait for Clk_period;
		Addr <=  "0001100011001";
		Trees_din <= x"ff790cc9";
		wait for Clk_period;
		Addr <=  "0001100011010";
		Trees_din <= x"001b0cc9";
		wait for Clk_period;
		Addr <=  "0001100011011";
		Trees_din <= x"a3ff8904";
		wait for Clk_period;
		Addr <=  "0001100011100";
		Trees_din <= x"ffc10cc9";
		wait for Clk_period;
		Addr <=  "0001100011101";
		Trees_din <= x"008a0cc9";
		wait for Clk_period;
		Addr <=  "0001100011110";
		Trees_din <= x"f9000d08";
		wait for Clk_period;
		Addr <=  "0001100011111";
		Trees_din <= x"f2037004";
		wait for Clk_period;
		Addr <=  "0001100100000";
		Trees_din <= x"ff6f0cc9";
		wait for Clk_period;
		Addr <=  "0001100100001";
		Trees_din <= x"00120cc9";
		wait for Clk_period;
		Addr <=  "0001100100010";
		Trees_din <= x"ddfe9a04";
		wait for Clk_period;
		Addr <=  "0001100100011";
		Trees_din <= x"01b70cc9";
		wait for Clk_period;
		Addr <=  "0001100100100";
		Trees_din <= x"ff9c0cc9";
		wait for Clk_period;
		Addr <=  "0001100100101";
		Trees_din <= x"37ff6d10";
		wait for Clk_period;
		Addr <=  "0001100100110";
		Trees_din <= x"fcfef008";
		wait for Clk_period;
		Addr <=  "0001100100111";
		Trees_din <= x"9fff7b04";
		wait for Clk_period;
		Addr <=  "0001100101000";
		Trees_din <= x"006b0cc9";
		wait for Clk_period;
		Addr <=  "0001100101001";
		Trees_din <= x"015e0cc9";
		wait for Clk_period;
		Addr <=  "0001100101010";
		Trees_din <= x"c8ffbc04";
		wait for Clk_period;
		Addr <=  "0001100101011";
		Trees_din <= x"009a0cc9";
		wait for Clk_period;
		Addr <=  "0001100101100";
		Trees_din <= x"ff7f0cc9";
		wait for Clk_period;
		Addr <=  "0001100101101";
		Trees_din <= x"3f008e08";
		wait for Clk_period;
		Addr <=  "0001100101110";
		Trees_din <= x"0dfeb604";
		wait for Clk_period;
		Addr <=  "0001100101111";
		Trees_din <= x"00650cc9";
		wait for Clk_period;
		Addr <=  "0001100110000";
		Trees_din <= x"ff7f0cc9";
		wait for Clk_period;
		Addr <=  "0001100110001";
		Trees_din <= x"00c90cc9";
		wait for Clk_period;
		Addr <=  "0001100110010";
		Trees_din <= x"00ff904c";
		wait for Clk_period;
		Addr <=  "0001100110011";
		Trees_din <= x"2f001a34";
		wait for Clk_period;
		Addr <=  "0001100110100";
		Trees_din <= x"8800ff20";
		wait for Clk_period;
		Addr <=  "0001100110101";
		Trees_din <= x"87ffcf10";
		wait for Clk_period;
		Addr <=  "0001100110110";
		Trees_din <= x"c6fe1108";
		wait for Clk_period;
		Addr <=  "0001100110111";
		Trees_din <= x"f3ff2d04";
		wait for Clk_period;
		Addr <=  "0001100111000";
		Trees_din <= x"ffad0e0d";
		wait for Clk_period;
		Addr <=  "0001100111001";
		Trees_din <= x"00dd0e0d";
		wait for Clk_period;
		Addr <=  "0001100111010";
		Trees_din <= x"ccff2c04";
		wait for Clk_period;
		Addr <=  "0001100111011";
		Trees_din <= x"fff20e0d";
		wait for Clk_period;
		Addr <=  "0001100111100";
		Trees_din <= x"ff830e0d";
		wait for Clk_period;
		Addr <=  "0001100111101";
		Trees_din <= x"74ffe108";
		wait for Clk_period;
		Addr <=  "0001100111110";
		Trees_din <= x"d6001904";
		wait for Clk_period;
		Addr <=  "0001100111111";
		Trees_din <= x"ffbb0e0d";
		wait for Clk_period;
		Addr <=  "0001101000000";
		Trees_din <= x"01140e0d";
		wait for Clk_period;
		Addr <=  "0001101000001";
		Trees_din <= x"3a000c04";
		wait for Clk_period;
		Addr <=  "0001101000010";
		Trees_din <= x"ff720e0d";
		wait for Clk_period;
		Addr <=  "0001101000011";
		Trees_din <= x"00430e0d";
		wait for Clk_period;
		Addr <=  "0001101000100";
		Trees_din <= x"e1ffe408";
		wait for Clk_period;
		Addr <=  "0001101000101";
		Trees_din <= x"10008d04";
		wait for Clk_period;
		Addr <=  "0001101000110";
		Trees_din <= x"ff860e0d";
		wait for Clk_period;
		Addr <=  "0001101000111";
		Trees_din <= x"00560e0d";
		wait for Clk_period;
		Addr <=  "0001101001000";
		Trees_din <= x"6e006708";
		wait for Clk_period;
		Addr <=  "0001101001001";
		Trees_din <= x"55ffce04";
		wait for Clk_period;
		Addr <=  "0001101001010";
		Trees_din <= x"00f80e0d";
		wait for Clk_period;
		Addr <=  "0001101001011";
		Trees_din <= x"00390e0d";
		wait for Clk_period;
		Addr <=  "0001101001100";
		Trees_din <= x"ffd90e0d";
		wait for Clk_period;
		Addr <=  "0001101001101";
		Trees_din <= x"7fff8f08";
		wait for Clk_period;
		Addr <=  "0001101001110";
		Trees_din <= x"9bffb804";
		wait for Clk_period;
		Addr <=  "0001101001111";
		Trees_din <= x"ff860e0d";
		wait for Clk_period;
		Addr <=  "0001101010000";
		Trees_din <= x"00450e0d";
		wait for Clk_period;
		Addr <=  "0001101010001";
		Trees_din <= x"f3fea404";
		wait for Clk_period;
		Addr <=  "0001101010010";
		Trees_din <= x"ffb00e0d";
		wait for Clk_period;
		Addr <=  "0001101010011";
		Trees_din <= x"68ff0e08";
		wait for Clk_period;
		Addr <=  "0001101010100";
		Trees_din <= x"28ff2a04";
		wait for Clk_period;
		Addr <=  "0001101010101";
		Trees_din <= x"003a0e0d";
		wait for Clk_period;
		Addr <=  "0001101010110";
		Trees_din <= x"01020e0d";
		wait for Clk_period;
		Addr <=  "0001101010111";
		Trees_din <= x"001d0e0d";
		wait for Clk_period;
		Addr <=  "0001101011000";
		Trees_din <= x"4bff102c";
		wait for Clk_period;
		Addr <=  "0001101011001";
		Trees_din <= x"65ff851c";
		wait for Clk_period;
		Addr <=  "0001101011010";
		Trees_din <= x"8dfe920c";
		wait for Clk_period;
		Addr <=  "0001101011011";
		Trees_din <= x"43fe8604";
		wait for Clk_period;
		Addr <=  "0001101011100";
		Trees_din <= x"00c80e0d";
		wait for Clk_period;
		Addr <=  "0001101011101";
		Trees_din <= x"e6ff7404";
		wait for Clk_period;
		Addr <=  "0001101011110";
		Trees_din <= x"00390e0d";
		wait for Clk_period;
		Addr <=  "0001101011111";
		Trees_din <= x"ff9a0e0d";
		wait for Clk_period;
		Addr <=  "0001101100000";
		Trees_din <= x"7bff8908";
		wait for Clk_period;
		Addr <=  "0001101100001";
		Trees_din <= x"c2fee304";
		wait for Clk_period;
		Addr <=  "0001101100010";
		Trees_din <= x"ffd60e0d";
		wait for Clk_period;
		Addr <=  "0001101100011";
		Trees_din <= x"00c00e0d";
		wait for Clk_period;
		Addr <=  "0001101100100";
		Trees_din <= x"51008004";
		wait for Clk_period;
		Addr <=  "0001101100101";
		Trees_din <= x"ff8d0e0d";
		wait for Clk_period;
		Addr <=  "0001101100110";
		Trees_din <= x"00600e0d";
		wait for Clk_period;
		Addr <=  "0001101100111";
		Trees_din <= x"86ffcb08";
		wait for Clk_period;
		Addr <=  "0001101101000";
		Trees_din <= x"00ff9304";
		wait for Clk_period;
		Addr <=  "0001101101001";
		Trees_din <= x"00760e0d";
		wait for Clk_period;
		Addr <=  "0001101101010";
		Trees_din <= x"ff6a0e0d";
		wait for Clk_period;
		Addr <=  "0001101101011";
		Trees_din <= x"14ff3404";
		wait for Clk_period;
		Addr <=  "0001101101100";
		Trees_din <= x"ffd40e0d";
		wait for Clk_period;
		Addr <=  "0001101101101";
		Trees_din <= x"00d30e0d";
		wait for Clk_period;
		Addr <=  "0001101101110";
		Trees_din <= x"90fffb14";
		wait for Clk_period;
		Addr <=  "0001101101111";
		Trees_din <= x"87fffa10";
		wait for Clk_period;
		Addr <=  "0001101110000";
		Trees_din <= x"fdffd108";
		wait for Clk_period;
		Addr <=  "0001101110001";
		Trees_din <= x"39feb704";
		wait for Clk_period;
		Addr <=  "0001101110010";
		Trees_din <= x"000f0e0d";
		wait for Clk_period;
		Addr <=  "0001101110011";
		Trees_din <= x"ff660e0d";
		wait for Clk_period;
		Addr <=  "0001101110100";
		Trees_din <= x"d8008904";
		wait for Clk_period;
		Addr <=  "0001101110101";
		Trees_din <= x"ff8b0e0d";
		wait for Clk_period;
		Addr <=  "0001101110110";
		Trees_din <= x"008b0e0d";
		wait for Clk_period;
		Addr <=  "0001101110111";
		Trees_din <= x"00850e0d";
		wait for Clk_period;
		Addr <=  "0001101111000";
		Trees_din <= x"b5ff0c10";
		wait for Clk_period;
		Addr <=  "0001101111001";
		Trees_din <= x"99ff1208";
		wait for Clk_period;
		Addr <=  "0001101111010";
		Trees_din <= x"74003204";
		wait for Clk_period;
		Addr <=  "0001101111011";
		Trees_din <= x"ffab0e0d";
		wait for Clk_period;
		Addr <=  "0001101111100";
		Trees_din <= x"00660e0d";
		wait for Clk_period;
		Addr <=  "0001101111101";
		Trees_din <= x"c6ff9c04";
		wait for Clk_period;
		Addr <=  "0001101111110";
		Trees_din <= x"00d60e0d";
		wait for Clk_period;
		Addr <=  "0001101111111";
		Trees_din <= x"fff70e0d";
		wait for Clk_period;
		Addr <=  "0001110000000";
		Trees_din <= x"6afedf04";
		wait for Clk_period;
		Addr <=  "0001110000001";
		Trees_din <= x"00430e0d";
		wait for Clk_period;
		Addr <=  "0001110000010";
		Trees_din <= x"ff750e0d";
		wait for Clk_period;
		Addr <=  "0001110000011";
		Trees_din <= x"00ff4140";
		wait for Clk_period;
		Addr <=  "0001110000100";
		Trees_din <= x"e1000a1c";
		wait for Clk_period;
		Addr <=  "0001110000101";
		Trees_din <= x"dc00ed14";
		wait for Clk_period;
		Addr <=  "0001110000110";
		Trees_din <= x"89010610";
		wait for Clk_period;
		Addr <=  "0001110000111";
		Trees_din <= x"bb003708";
		wait for Clk_period;
		Addr <=  "0001110001000";
		Trees_din <= x"ab015504";
		wait for Clk_period;
		Addr <=  "0001110001001";
		Trees_din <= x"ff660f79";
		wait for Clk_period;
		Addr <=  "0001110001010";
		Trees_din <= x"00170f79";
		wait for Clk_period;
		Addr <=  "0001110001011";
		Trees_din <= x"05ffeb04";
		wait for Clk_period;
		Addr <=  "0001110001100";
		Trees_din <= x"008d0f79";
		wait for Clk_period;
		Addr <=  "0001110001101";
		Trees_din <= x"ffa20f79";
		wait for Clk_period;
		Addr <=  "0001110001110";
		Trees_din <= x"00380f79";
		wait for Clk_period;
		Addr <=  "0001110001111";
		Trees_din <= x"e4fef704";
		wait for Clk_period;
		Addr <=  "0001110010000";
		Trees_din <= x"ffcd0f79";
		wait for Clk_period;
		Addr <=  "0001110010001";
		Trees_din <= x"009b0f79";
		wait for Clk_period;
		Addr <=  "0001110010010";
		Trees_din <= x"1f002f10";
		wait for Clk_period;
		Addr <=  "0001110010011";
		Trees_din <= x"e2fea508";
		wait for Clk_period;
		Addr <=  "0001110010100";
		Trees_din <= x"9dffc204";
		wait for Clk_period;
		Addr <=  "0001110010101";
		Trees_din <= x"ffa70f79";
		wait for Clk_period;
		Addr <=  "0001110010110";
		Trees_din <= x"00980f79";
		wait for Clk_period;
		Addr <=  "0001110010111";
		Trees_din <= x"8aff2104";
		wait for Clk_period;
		Addr <=  "0001110011000";
		Trees_din <= x"ffed0f79";
		wait for Clk_period;
		Addr <=  "0001110011001";
		Trees_din <= x"ff720f79";
		wait for Clk_period;
		Addr <=  "0001110011010";
		Trees_din <= x"2affca0c";
		wait for Clk_period;
		Addr <=  "0001110011011";
		Trees_din <= x"76ffa408";
		wait for Clk_period;
		Addr <=  "0001110011100";
		Trees_din <= x"03003604";
		wait for Clk_period;
		Addr <=  "0001110011101";
		Trees_din <= x"01d60f79";
		wait for Clk_period;
		Addr <=  "0001110011110";
		Trees_din <= x"00890f79";
		wait for Clk_period;
		Addr <=  "0001110011111";
		Trees_din <= x"fff00f79";
		wait for Clk_period;
		Addr <=  "0001110100000";
		Trees_din <= x"c3ff5904";
		wait for Clk_period;
		Addr <=  "0001110100001";
		Trees_din <= x"008a0f79";
		wait for Clk_period;
		Addr <=  "0001110100010";
		Trees_din <= x"ff870f79";
		wait for Clk_period;
		Addr <=  "0001110100011";
		Trees_din <= x"c7fee63c";
		wait for Clk_period;
		Addr <=  "0001110100100";
		Trees_din <= x"8dfe641c";
		wait for Clk_period;
		Addr <=  "0001110100101";
		Trees_din <= x"e6ff9d10";
		wait for Clk_period;
		Addr <=  "0001110100110";
		Trees_din <= x"89004208";
		wait for Clk_period;
		Addr <=  "0001110100111";
		Trees_din <= x"04ff9204";
		wait for Clk_period;
		Addr <=  "0001110101000";
		Trees_din <= x"00bd0f79";
		wait for Clk_period;
		Addr <=  "0001110101001";
		Trees_din <= x"ff720f79";
		wait for Clk_period;
		Addr <=  "0001110101010";
		Trees_din <= x"95ff2d04";
		wait for Clk_period;
		Addr <=  "0001110101011";
		Trees_din <= x"ffdc0f79";
		wait for Clk_period;
		Addr <=  "0001110101100";
		Trees_din <= x"009c0f79";
		wait for Clk_period;
		Addr <=  "0001110101101";
		Trees_din <= x"69fe4b04";
		wait for Clk_period;
		Addr <=  "0001110101110";
		Trees_din <= x"00690f79";
		wait for Clk_period;
		Addr <=  "0001110101111";
		Trees_din <= x"90fffb04";
		wait for Clk_period;
		Addr <=  "0001110110000";
		Trees_din <= x"ff6b0f79";
		wait for Clk_period;
		Addr <=  "0001110110001";
		Trees_din <= x"ffde0f79";
		wait for Clk_period;
		Addr <=  "0001110110010";
		Trees_din <= x"43ff6c10";
		wait for Clk_period;
		Addr <=  "0001110110011";
		Trees_din <= x"90ff6208";
		wait for Clk_period;
		Addr <=  "0001110110100";
		Trees_din <= x"2f000504";
		wait for Clk_period;
		Addr <=  "0001110110101";
		Trees_din <= x"ff760f79";
		wait for Clk_period;
		Addr <=  "0001110110110";
		Trees_din <= x"002a0f79";
		wait for Clk_period;
		Addr <=  "0001110110111";
		Trees_din <= x"2eff6d04";
		wait for Clk_period;
		Addr <=  "0001110111000";
		Trees_din <= x"ff7d0f79";
		wait for Clk_period;
		Addr <=  "0001110111001";
		Trees_din <= x"00580f79";
		wait for Clk_period;
		Addr <=  "0001110111010";
		Trees_din <= x"f800b708";
		wait for Clk_period;
		Addr <=  "0001110111011";
		Trees_din <= x"2cffcc04";
		wait for Clk_period;
		Addr <=  "0001110111100";
		Trees_din <= x"00130f79";
		wait for Clk_period;
		Addr <=  "0001110111101";
		Trees_din <= x"00ad0f79";
		wait for Clk_period;
		Addr <=  "0001110111110";
		Trees_din <= x"1dfec604";
		wait for Clk_period;
		Addr <=  "0001110111111";
		Trees_din <= x"02030f79";
		wait for Clk_period;
		Addr <=  "0001111000000";
		Trees_din <= x"00790f79";
		wait for Clk_period;
		Addr <=  "0001111000001";
		Trees_din <= x"51007020";
		wait for Clk_period;
		Addr <=  "0001111000010";
		Trees_din <= x"c6feb510";
		wait for Clk_period;
		Addr <=  "0001111000011";
		Trees_din <= x"cdffdd08";
		wait for Clk_period;
		Addr <=  "0001111000100";
		Trees_din <= x"79fec204";
		wait for Clk_period;
		Addr <=  "0001111000101";
		Trees_din <= x"00340f79";
		wait for Clk_period;
		Addr <=  "0001111000110";
		Trees_din <= x"ff8a0f79";
		wait for Clk_period;
		Addr <=  "0001111000111";
		Trees_din <= x"1cff3704";
		wait for Clk_period;
		Addr <=  "0001111001000";
		Trees_din <= x"01000f79";
		wait for Clk_period;
		Addr <=  "0001111001001";
		Trees_din <= x"00070f79";
		wait for Clk_period;
		Addr <=  "0001111001010";
		Trees_din <= x"b0fec708";
		wait for Clk_period;
		Addr <=  "0001111001011";
		Trees_din <= x"d000e704";
		wait for Clk_period;
		Addr <=  "0001111001100";
		Trees_din <= x"ffab0f79";
		wait for Clk_period;
		Addr <=  "0001111001101";
		Trees_din <= x"00b10f79";
		wait for Clk_period;
		Addr <=  "0001111001110";
		Trees_din <= x"f2036704";
		wait for Clk_period;
		Addr <=  "0001111001111";
		Trees_din <= x"ff800f79";
		wait for Clk_period;
		Addr <=  "0001111010000";
		Trees_din <= x"00470f79";
		wait for Clk_period;
		Addr <=  "0001111010001";
		Trees_din <= x"7fffb310";
		wait for Clk_period;
		Addr <=  "0001111010010";
		Trees_din <= x"71ff1f08";
		wait for Clk_period;
		Addr <=  "0001111010011";
		Trees_din <= x"43ffb904";
		wait for Clk_period;
		Addr <=  "0001111010100";
		Trees_din <= x"ffb40f79";
		wait for Clk_period;
		Addr <=  "0001111010101";
		Trees_din <= x"00a40f79";
		wait for Clk_period;
		Addr <=  "0001111010110";
		Trees_din <= x"d3ff5504";
		wait for Clk_period;
		Addr <=  "0001111010111";
		Trees_din <= x"ff780f79";
		wait for Clk_period;
		Addr <=  "0001111011000";
		Trees_din <= x"fffe0f79";
		wait for Clk_period;
		Addr <=  "0001111011001";
		Trees_din <= x"aaff4e04";
		wait for Clk_period;
		Addr <=  "0001111011010";
		Trees_din <= x"ff9c0f79";
		wait for Clk_period;
		Addr <=  "0001111011011";
		Trees_din <= x"66ffab04";
		wait for Clk_period;
		Addr <=  "0001111011100";
		Trees_din <= x"001a0f79";
		wait for Clk_period;
		Addr <=  "0001111011101";
		Trees_din <= x"00f40f79";
		wait for Clk_period;
		Addr <=  "0001111011110";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0001111011111";
		Trees_din <= x"00ff4138";
		wait for Clk_period;
		Addr <=  "0001111100000";
		Trees_din <= x"e1000a1c";
		wait for Clk_period;
		Addr <=  "0001111100001";
		Trees_din <= x"dc00ed14";
		wait for Clk_period;
		Addr <=  "0001111100010";
		Trees_din <= x"89010610";
		wait for Clk_period;
		Addr <=  "0001111100011";
		Trees_din <= x"dffeec08";
		wait for Clk_period;
		Addr <=  "0001111100100";
		Trees_din <= x"51005004";
		wait for Clk_period;
		Addr <=  "0001111100101";
		Trees_din <= x"ff8810c1";
		wait for Clk_period;
		Addr <=  "0001111100110";
		Trees_din <= x"009510c1";
		wait for Clk_period;
		Addr <=  "0001111100111";
		Trees_din <= x"b4fdb404";
		wait for Clk_period;
		Addr <=  "0001111101000";
		Trees_din <= x"fff710c1";
		wait for Clk_period;
		Addr <=  "0001111101001";
		Trees_din <= x"ff6610c1";
		wait for Clk_period;
		Addr <=  "0001111101010";
		Trees_din <= x"003410c1";
		wait for Clk_period;
		Addr <=  "0001111101011";
		Trees_din <= x"e4fef704";
		wait for Clk_period;
		Addr <=  "0001111101100";
		Trees_din <= x"ffd110c1";
		wait for Clk_period;
		Addr <=  "0001111101101";
		Trees_din <= x"008b10c1";
		wait for Clk_period;
		Addr <=  "0001111101110";
		Trees_din <= x"1f002f0c";
		wait for Clk_period;
		Addr <=  "0001111101111";
		Trees_din <= x"a7feb204";
		wait for Clk_period;
		Addr <=  "0001111110000";
		Trees_din <= x"008510c1";
		wait for Clk_period;
		Addr <=  "0001111110001";
		Trees_din <= x"1afe4d04";
		wait for Clk_period;
		Addr <=  "0001111110010";
		Trees_din <= x"002a10c1";
		wait for Clk_period;
		Addr <=  "0001111110011";
		Trees_din <= x"ff7310c1";
		wait for Clk_period;
		Addr <=  "0001111110100";
		Trees_din <= x"9cff9204";
		wait for Clk_period;
		Addr <=  "0001111110101";
		Trees_din <= x"ff9410c1";
		wait for Clk_period;
		Addr <=  "0001111110110";
		Trees_din <= x"b7ff8b04";
		wait for Clk_period;
		Addr <=  "0001111110111";
		Trees_din <= x"ffe010c1";
		wait for Clk_period;
		Addr <=  "0001111111000";
		Trees_din <= x"76ffa404";
		wait for Clk_period;
		Addr <=  "0001111111001";
		Trees_din <= x"014f10c1";
		wait for Clk_period;
		Addr <=  "0001111111010";
		Trees_din <= x"003b10c1";
		wait for Clk_period;
		Addr <=  "0001111111011";
		Trees_din <= x"c7fee634";
		wait for Clk_period;
		Addr <=  "0001111111100";
		Trees_din <= x"43ffa920";
		wait for Clk_period;
		Addr <=  "0001111111101";
		Trees_din <= x"5cff9c10";
		wait for Clk_period;
		Addr <=  "0001111111110";
		Trees_din <= x"37ff7608";
		wait for Clk_period;
		Addr <=  "0001111111111";
		Trees_din <= x"ebfeb904";
		wait for Clk_period;
		Addr <=  "0010000000000";
		Trees_din <= x"ffc310c1";
		wait for Clk_period;
		Addr <=  "0010000000001";
		Trees_din <= x"00d810c1";
		wait for Clk_period;
		Addr <=  "0010000000010";
		Trees_din <= x"dc00ed04";
		wait for Clk_period;
		Addr <=  "0010000000011";
		Trees_din <= x"ff8210c1";
		wait for Clk_period;
		Addr <=  "0010000000100";
		Trees_din <= x"007810c1";
		wait for Clk_period;
		Addr <=  "0010000000101";
		Trees_din <= x"ccff3f08";
		wait for Clk_period;
		Addr <=  "0010000000110";
		Trees_din <= x"54005804";
		wait for Clk_period;
		Addr <=  "0010000000111";
		Trees_din <= x"ffc710c1";
		wait for Clk_period;
		Addr <=  "0010000001000";
		Trees_din <= x"009a10c1";
		wait for Clk_period;
		Addr <=  "0010000001001";
		Trees_din <= x"d000c204";
		wait for Clk_period;
		Addr <=  "0010000001010";
		Trees_din <= x"ff6f10c1";
		wait for Clk_period;
		Addr <=  "0010000001011";
		Trees_din <= x"000010c1";
		wait for Clk_period;
		Addr <=  "0010000001100";
		Trees_din <= x"59001910";
		wait for Clk_period;
		Addr <=  "0010000001101";
		Trees_din <= x"14ff3d08";
		wait for Clk_period;
		Addr <=  "0010000001110";
		Trees_din <= x"79fed104";
		wait for Clk_period;
		Addr <=  "0010000001111";
		Trees_din <= x"000710c1";
		wait for Clk_period;
		Addr <=  "0010000010000";
		Trees_din <= x"00b710c1";
		wait for Clk_period;
		Addr <=  "0010000010001";
		Trees_din <= x"5e000404";
		wait for Clk_period;
		Addr <=  "0010000010010";
		Trees_din <= x"ff8c10c1";
		wait for Clk_period;
		Addr <=  "0010000010011";
		Trees_din <= x"006a10c1";
		wait for Clk_period;
		Addr <=  "0010000010100";
		Trees_din <= x"ff8c10c1";
		wait for Clk_period;
		Addr <=  "0010000010101";
		Trees_din <= x"1afeca20";
		wait for Clk_period;
		Addr <=  "0010000010110";
		Trees_din <= x"88001110";
		wait for Clk_period;
		Addr <=  "0010000010111";
		Trees_din <= x"60ff0808";
		wait for Clk_period;
		Addr <=  "0010000011000";
		Trees_din <= x"dcff5804";
		wait for Clk_period;
		Addr <=  "0010000011001";
		Trees_din <= x"010f10c1";
		wait for Clk_period;
		Addr <=  "0010000011010";
		Trees_din <= x"ffae10c1";
		wait for Clk_period;
		Addr <=  "0010000011011";
		Trees_din <= x"51009104";
		wait for Clk_period;
		Addr <=  "0010000011100";
		Trees_din <= x"ff6e10c1";
		wait for Clk_period;
		Addr <=  "0010000011101";
		Trees_din <= x"001910c1";
		wait for Clk_period;
		Addr <=  "0010000011110";
		Trees_din <= x"e9ff2508";
		wait for Clk_period;
		Addr <=  "0010000011111";
		Trees_din <= x"c0ff5804";
		wait for Clk_period;
		Addr <=  "0010000100000";
		Trees_din <= x"000810c1";
		wait for Clk_period;
		Addr <=  "0010000100001";
		Trees_din <= x"00b610c1";
		wait for Clk_period;
		Addr <=  "0010000100010";
		Trees_din <= x"f6feb404";
		wait for Clk_period;
		Addr <=  "0010000100011";
		Trees_din <= x"006710c1";
		wait for Clk_period;
		Addr <=  "0010000100100";
		Trees_din <= x"ff8210c1";
		wait for Clk_period;
		Addr <=  "0010000100101";
		Trees_din <= x"c6fead0c";
		wait for Clk_period;
		Addr <=  "0010000100110";
		Trees_din <= x"ac004504";
		wait for Clk_period;
		Addr <=  "0010000100111";
		Trees_din <= x"ffcb10c1";
		wait for Clk_period;
		Addr <=  "0010000101000";
		Trees_din <= x"daffc404";
		wait for Clk_period;
		Addr <=  "0010000101001";
		Trees_din <= x"010610c1";
		wait for Clk_period;
		Addr <=  "0010000101010";
		Trees_din <= x"003110c1";
		wait for Clk_period;
		Addr <=  "0010000101011";
		Trees_din <= x"1200bd08";
		wait for Clk_period;
		Addr <=  "0010000101100";
		Trees_din <= x"5affab04";
		wait for Clk_period;
		Addr <=  "0010000101101";
		Trees_din <= x"001d10c1";
		wait for Clk_period;
		Addr <=  "0010000101110";
		Trees_din <= x"ff6f10c1";
		wait for Clk_period;
		Addr <=  "0010000101111";
		Trees_din <= x"005710c1";
		wait for Clk_period;
		Addr <=  "0010000110000";
		Trees_din <= x"0fff3148";
		wait for Clk_period;
		Addr <=  "0010000110001";
		Trees_din <= x"1cfee118";
		wait for Clk_period;
		Addr <=  "0010000110010";
		Trees_din <= x"aaff0904";
		wait for Clk_period;
		Addr <=  "0010000110011";
		Trees_din <= x"ffae11fd";
		wait for Clk_period;
		Addr <=  "0010000110100";
		Trees_din <= x"d8006510";
		wait for Clk_period;
		Addr <=  "0010000110101";
		Trees_din <= x"78ff5208";
		wait for Clk_period;
		Addr <=  "0010000110110";
		Trees_din <= x"7efe8104";
		wait for Clk_period;
		Addr <=  "0010000110111";
		Trees_din <= x"002f11fd";
		wait for Clk_period;
		Addr <=  "0010000111000";
		Trees_din <= x"00f311fd";
		wait for Clk_period;
		Addr <=  "0010000111001";
		Trees_din <= x"5a003904";
		wait for Clk_period;
		Addr <=  "0010000111010";
		Trees_din <= x"009511fd";
		wait for Clk_period;
		Addr <=  "0010000111011";
		Trees_din <= x"ffab11fd";
		wait for Clk_period;
		Addr <=  "0010000111100";
		Trees_din <= x"ffee11fd";
		wait for Clk_period;
		Addr <=  "0010000111101";
		Trees_din <= x"07002d10";
		wait for Clk_period;
		Addr <=  "0010000111110";
		Trees_din <= x"4dfdfc04";
		wait for Clk_period;
		Addr <=  "0010000111111";
		Trees_din <= x"009211fd";
		wait for Clk_period;
		Addr <=  "0010001000000";
		Trees_din <= x"3bfe7204";
		wait for Clk_period;
		Addr <=  "0010001000001";
		Trees_din <= x"004711fd";
		wait for Clk_period;
		Addr <=  "0010001000010";
		Trees_din <= x"39fef704";
		wait for Clk_period;
		Addr <=  "0010001000011";
		Trees_din <= x"fff011fd";
		wait for Clk_period;
		Addr <=  "0010001000100";
		Trees_din <= x"ff6c11fd";
		wait for Clk_period;
		Addr <=  "0010001000101";
		Trees_din <= x"90ffad10";
		wait for Clk_period;
		Addr <=  "0010001000110";
		Trees_din <= x"f3ff2008";
		wait for Clk_period;
		Addr <=  "0010001000111";
		Trees_din <= x"ecff7904";
		wait for Clk_period;
		Addr <=  "0010001001000";
		Trees_din <= x"002a11fd";
		wait for Clk_period;
		Addr <=  "0010001001001";
		Trees_din <= x"ff7111fd";
		wait for Clk_period;
		Addr <=  "0010001001010";
		Trees_din <= x"ccff7104";
		wait for Clk_period;
		Addr <=  "0010001001011";
		Trees_din <= x"00aa11fd";
		wait for Clk_period;
		Addr <=  "0010001001100";
		Trees_din <= x"ffc611fd";
		wait for Clk_period;
		Addr <=  "0010001001101";
		Trees_din <= x"aeff2508";
		wait for Clk_period;
		Addr <=  "0010001001110";
		Trees_din <= x"8aff8b04";
		wait for Clk_period;
		Addr <=  "0010001001111";
		Trees_din <= x"ffe711fd";
		wait for Clk_period;
		Addr <=  "0010001010000";
		Trees_din <= x"009b11fd";
		wait for Clk_period;
		Addr <=  "0010001010001";
		Trees_din <= x"8e00bf04";
		wait for Clk_period;
		Addr <=  "0010001010010";
		Trees_din <= x"ffaa11fd";
		wait for Clk_period;
		Addr <=  "0010001010011";
		Trees_din <= x"005111fd";
		wait for Clk_period;
		Addr <=  "0010001010100";
		Trees_din <= x"30ffb51c";
		wait for Clk_period;
		Addr <=  "0010001010101";
		Trees_din <= x"2c006814";
		wait for Clk_period;
		Addr <=  "0010001010110";
		Trees_din <= x"90fea308";
		wait for Clk_period;
		Addr <=  "0010001010111";
		Trees_din <= x"b2005a04";
		wait for Clk_period;
		Addr <=  "0010001011000";
		Trees_din <= x"ff9d11fd";
		wait for Clk_period;
		Addr <=  "0010001011001";
		Trees_din <= x"009911fd";
		wait for Clk_period;
		Addr <=  "0010001011010";
		Trees_din <= x"35001608";
		wait for Clk_period;
		Addr <=  "0010001011011";
		Trees_din <= x"f8ff6204";
		wait for Clk_period;
		Addr <=  "0010001011100";
		Trees_din <= x"ffde11fd";
		wait for Clk_period;
		Addr <=  "0010001011101";
		Trees_din <= x"ff6611fd";
		wait for Clk_period;
		Addr <=  "0010001011110";
		Trees_din <= x"002a11fd";
		wait for Clk_period;
		Addr <=  "0010001011111";
		Trees_din <= x"50ff1f04";
		wait for Clk_period;
		Addr <=  "0010001100000";
		Trees_din <= x"00b111fd";
		wait for Clk_period;
		Addr <=  "0010001100001";
		Trees_din <= x"ffa211fd";
		wait for Clk_period;
		Addr <=  "0010001100010";
		Trees_din <= x"73ffd31c";
		wait for Clk_period;
		Addr <=  "0010001100011";
		Trees_din <= x"59ff4310";
		wait for Clk_period;
		Addr <=  "0010001100100";
		Trees_din <= x"51002b08";
		wait for Clk_period;
		Addr <=  "0010001100101";
		Trees_din <= x"e9ffe704";
		wait for Clk_period;
		Addr <=  "0010001100110";
		Trees_din <= x"ff7911fd";
		wait for Clk_period;
		Addr <=  "0010001100111";
		Trees_din <= x"006f11fd";
		wait for Clk_period;
		Addr <=  "0010001101000";
		Trees_din <= x"12ff8604";
		wait for Clk_period;
		Addr <=  "0010001101001";
		Trees_din <= x"00ef11fd";
		wait for Clk_period;
		Addr <=  "0010001101010";
		Trees_din <= x"ffc511fd";
		wait for Clk_period;
		Addr <=  "0010001101011";
		Trees_din <= x"10feb304";
		wait for Clk_period;
		Addr <=  "0010001101100";
		Trees_din <= x"005f11fd";
		wait for Clk_period;
		Addr <=  "0010001101101";
		Trees_din <= x"faffbe04";
		wait for Clk_period;
		Addr <=  "0010001101110";
		Trees_din <= x"ff6811fd";
		wait for Clk_period;
		Addr <=  "0010001101111";
		Trees_din <= x"ffdf11fd";
		wait for Clk_period;
		Addr <=  "0010001110000";
		Trees_din <= x"ac003710";
		wait for Clk_period;
		Addr <=  "0010001110001";
		Trees_din <= x"64ff2b08";
		wait for Clk_period;
		Addr <=  "0010001110010";
		Trees_din <= x"6d006204";
		wait for Clk_period;
		Addr <=  "0010001110011";
		Trees_din <= x"ffcb11fd";
		wait for Clk_period;
		Addr <=  "0010001110100";
		Trees_din <= x"009c11fd";
		wait for Clk_period;
		Addr <=  "0010001110101";
		Trees_din <= x"de00ad04";
		wait for Clk_period;
		Addr <=  "0010001110110";
		Trees_din <= x"ff6e11fd";
		wait for Clk_period;
		Addr <=  "0010001110111";
		Trees_din <= x"ffe511fd";
		wait for Clk_period;
		Addr <=  "0010001111000";
		Trees_din <= x"1eff9208";
		wait for Clk_period;
		Addr <=  "0010001111001";
		Trees_din <= x"a3002504";
		wait for Clk_period;
		Addr <=  "0010001111010";
		Trees_din <= x"ffb211fd";
		wait for Clk_period;
		Addr <=  "0010001111011";
		Trees_din <= x"00a211fd";
		wait for Clk_period;
		Addr <=  "0010001111100";
		Trees_din <= x"2affee04";
		wait for Clk_period;
		Addr <=  "0010001111101";
		Trees_din <= x"fff211fd";
		wait for Clk_period;
		Addr <=  "0010001111110";
		Trees_din <= x"00b611fd";
		wait for Clk_period;
		Addr <=  "0010001111111";
		Trees_din <= x"00ff4130";
		wait for Clk_period;
		Addr <=  "0010010000000";
		Trees_din <= x"e1000a18";
		wait for Clk_period;
		Addr <=  "0010010000001";
		Trees_din <= x"dc00ed10";
		wait for Clk_period;
		Addr <=  "0010010000010";
		Trees_din <= x"8901060c";
		wait for Clk_period;
		Addr <=  "0010010000011";
		Trees_din <= x"bb003708";
		wait for Clk_period;
		Addr <=  "0010010000100";
		Trees_din <= x"ab015504";
		wait for Clk_period;
		Addr <=  "0010010000101";
		Trees_din <= x"ff691301";
		wait for Clk_period;
		Addr <=  "0010010000110";
		Trees_din <= x"00141301";
		wait for Clk_period;
		Addr <=  "0010010000111";
		Trees_din <= x"00141301";
		wait for Clk_period;
		Addr <=  "0010010001000";
		Trees_din <= x"002f1301";
		wait for Clk_period;
		Addr <=  "0010010001001";
		Trees_din <= x"baff9004";
		wait for Clk_period;
		Addr <=  "0010010001010";
		Trees_din <= x"00701301";
		wait for Clk_period;
		Addr <=  "0010010001011";
		Trees_din <= x"ffe81301";
		wait for Clk_period;
		Addr <=  "0010010001100";
		Trees_din <= x"76ffa810";
		wait for Clk_period;
		Addr <=  "0010010001101";
		Trees_din <= x"1cff680c";
		wait for Clk_period;
		Addr <=  "0010010001110";
		Trees_din <= x"ccffb808";
		wait for Clk_period;
		Addr <=  "0010010001111";
		Trees_din <= x"5effac04";
		wait for Clk_period;
		Addr <=  "0010010010000";
		Trees_din <= x"000f1301";
		wait for Clk_period;
		Addr <=  "0010010010001";
		Trees_din <= x"00f01301";
		wait for Clk_period;
		Addr <=  "0010010010010";
		Trees_din <= x"ffe51301";
		wait for Clk_period;
		Addr <=  "0010010010011";
		Trees_din <= x"ff941301";
		wait for Clk_period;
		Addr <=  "0010010010100";
		Trees_din <= x"0b00bf04";
		wait for Clk_period;
		Addr <=  "0010010010101";
		Trees_din <= x"ff781301";
		wait for Clk_period;
		Addr <=  "0010010010110";
		Trees_din <= x"00621301";
		wait for Clk_period;
		Addr <=  "0010010010111";
		Trees_din <= x"c7ff0b24";
		wait for Clk_period;
		Addr <=  "0010010011000";
		Trees_din <= x"5900271c";
		wait for Clk_period;
		Addr <=  "0010010011001";
		Trees_din <= x"43ffa910";
		wait for Clk_period;
		Addr <=  "0010010011010";
		Trees_din <= x"7fffe608";
		wait for Clk_period;
		Addr <=  "0010010011011";
		Trees_din <= x"a3ff8504";
		wait for Clk_period;
		Addr <=  "0010010011100";
		Trees_din <= x"ffa51301";
		wait for Clk_period;
		Addr <=  "0010010011101";
		Trees_din <= x"00211301";
		wait for Clk_period;
		Addr <=  "0010010011110";
		Trees_din <= x"c5ff3104";
		wait for Clk_period;
		Addr <=  "0010010011111";
		Trees_din <= x"00c01301";
		wait for Clk_period;
		Addr <=  "0010010100000";
		Trees_din <= x"ffd61301";
		wait for Clk_period;
		Addr <=  "0010010100001";
		Trees_din <= x"0fffee08";
		wait for Clk_period;
		Addr <=  "0010010100010";
		Trees_din <= x"f4fed604";
		wait for Clk_period;
		Addr <=  "0010010100011";
		Trees_din <= x"00a61301";
		wait for Clk_period;
		Addr <=  "0010010100100";
		Trees_din <= x"00401301";
		wait for Clk_period;
		Addr <=  "0010010100101";
		Trees_din <= x"ffa01301";
		wait for Clk_period;
		Addr <=  "0010010100110";
		Trees_din <= x"43fe7b04";
		wait for Clk_period;
		Addr <=  "0010010100111";
		Trees_din <= x"00561301";
		wait for Clk_period;
		Addr <=  "0010010101000";
		Trees_din <= x"ff701301";
		wait for Clk_period;
		Addr <=  "0010010101001";
		Trees_din <= x"9cff9618";
		wait for Clk_period;
		Addr <=  "0010010101010";
		Trees_din <= x"50fef00c";
		wait for Clk_period;
		Addr <=  "0010010101011";
		Trees_din <= x"68fe4f04";
		wait for Clk_period;
		Addr <=  "0010010101100";
		Trees_din <= x"00bc1301";
		wait for Clk_period;
		Addr <=  "0010010101101";
		Trees_din <= x"89008a04";
		wait for Clk_period;
		Addr <=  "0010010101110";
		Trees_din <= x"ff8f1301";
		wait for Clk_period;
		Addr <=  "0010010101111";
		Trees_din <= x"002d1301";
		wait for Clk_period;
		Addr <=  "0010010110000";
		Trees_din <= x"d9003e08";
		wait for Clk_period;
		Addr <=  "0010010110001";
		Trees_din <= x"70fde604";
		wait for Clk_period;
		Addr <=  "0010010110010";
		Trees_din <= x"00111301";
		wait for Clk_period;
		Addr <=  "0010010110011";
		Trees_din <= x"ff701301";
		wait for Clk_period;
		Addr <=  "0010010110100";
		Trees_din <= x"004d1301";
		wait for Clk_period;
		Addr <=  "0010010110101";
		Trees_din <= x"c3ffe310";
		wait for Clk_period;
		Addr <=  "0010010110110";
		Trees_din <= x"f7ff9b08";
		wait for Clk_period;
		Addr <=  "0010010110111";
		Trees_din <= x"aaff7204";
		wait for Clk_period;
		Addr <=  "0010010111000";
		Trees_din <= x"ffdb1301";
		wait for Clk_period;
		Addr <=  "0010010111001";
		Trees_din <= x"00b31301";
		wait for Clk_period;
		Addr <=  "0010010111010";
		Trees_din <= x"65ff1104";
		wait for Clk_period;
		Addr <=  "0010010111011";
		Trees_din <= x"003e1301";
		wait for Clk_period;
		Addr <=  "0010010111100";
		Trees_din <= x"ff821301";
		wait for Clk_period;
		Addr <=  "0010010111101";
		Trees_din <= x"b8002504";
		wait for Clk_period;
		Addr <=  "0010010111110";
		Trees_din <= x"ff721301";
		wait for Clk_period;
		Addr <=  "0010010111111";
		Trees_din <= x"00911301";
		wait for Clk_period;
		Addr <=  "0010011000000";
		Trees_din <= x"0dff6958";
		wait for Clk_period;
		Addr <=  "0010011000001";
		Trees_din <= x"30ffb520";
		wait for Clk_period;
		Addr <=  "0010011000010";
		Trees_din <= x"0fff2b14";
		wait for Clk_period;
		Addr <=  "0010011000011";
		Trees_din <= x"b9feda0c";
		wait for Clk_period;
		Addr <=  "0010011000100";
		Trees_din <= x"e4fe9908";
		wait for Clk_period;
		Addr <=  "0010011000101";
		Trees_din <= x"daffdf04";
		wait for Clk_period;
		Addr <=  "0010011000110";
		Trees_din <= x"ffea1445";
		wait for Clk_period;
		Addr <=  "0010011000111";
		Trees_din <= x"00af1445";
		wait for Clk_period;
		Addr <=  "0010011001000";
		Trees_din <= x"ffdf1445";
		wait for Clk_period;
		Addr <=  "0010011001001";
		Trees_din <= x"ceff1404";
		wait for Clk_period;
		Addr <=  "0010011001010";
		Trees_din <= x"004a1445";
		wait for Clk_period;
		Addr <=  "0010011001011";
		Trees_din <= x"ff831445";
		wait for Clk_period;
		Addr <=  "0010011001100";
		Trees_din <= x"3d00a608";
		wait for Clk_period;
		Addr <=  "0010011001101";
		Trees_din <= x"2c006804";
		wait for Clk_period;
		Addr <=  "0010011001110";
		Trees_din <= x"ff6b1445";
		wait for Clk_period;
		Addr <=  "0010011001111";
		Trees_din <= x"00111445";
		wait for Clk_period;
		Addr <=  "0010011010000";
		Trees_din <= x"00681445";
		wait for Clk_period;
		Addr <=  "0010011010001";
		Trees_din <= x"87ff9a20";
		wait for Clk_period;
		Addr <=  "0010011010010";
		Trees_din <= x"88006c10";
		wait for Clk_period;
		Addr <=  "0010011010011";
		Trees_din <= x"b4fe8908";
		wait for Clk_period;
		Addr <=  "0010011010100";
		Trees_din <= x"64fec004";
		wait for Clk_period;
		Addr <=  "0010011010101";
		Trees_din <= x"00931445";
		wait for Clk_period;
		Addr <=  "0010011010110";
		Trees_din <= x"fff41445";
		wait for Clk_period;
		Addr <=  "0010011010111";
		Trees_din <= x"36fef104";
		wait for Clk_period;
		Addr <=  "0010011011000";
		Trees_din <= x"00191445";
		wait for Clk_period;
		Addr <=  "0010011011001";
		Trees_din <= x"ff8e1445";
		wait for Clk_period;
		Addr <=  "0010011011010";
		Trees_din <= x"6affb008";
		wait for Clk_period;
		Addr <=  "0010011011011";
		Trees_din <= x"68fe9704";
		wait for Clk_period;
		Addr <=  "0010011011100";
		Trees_din <= x"00b91445";
		wait for Clk_period;
		Addr <=  "0010011011101";
		Trees_din <= x"003b1445";
		wait for Clk_period;
		Addr <=  "0010011011110";
		Trees_din <= x"a7ffeb04";
		wait for Clk_period;
		Addr <=  "0010011011111";
		Trees_din <= x"ff841445";
		wait for Clk_period;
		Addr <=  "0010011100000";
		Trees_din <= x"00351445";
		wait for Clk_period;
		Addr <=  "0010011100001";
		Trees_din <= x"adff3e08";
		wait for Clk_period;
		Addr <=  "0010011100010";
		Trees_din <= x"c8005004";
		wait for Clk_period;
		Addr <=  "0010011100011";
		Trees_din <= x"ff8d1445";
		wait for Clk_period;
		Addr <=  "0010011100100";
		Trees_din <= x"00491445";
		wait for Clk_period;
		Addr <=  "0010011100101";
		Trees_din <= x"2affca08";
		wait for Clk_period;
		Addr <=  "0010011100110";
		Trees_din <= x"a6ff8704";
		wait for Clk_period;
		Addr <=  "0010011100111";
		Trees_din <= x"ff9e1445";
		wait for Clk_period;
		Addr <=  "0010011101000";
		Trees_din <= x"005e1445";
		wait for Clk_period;
		Addr <=  "0010011101001";
		Trees_din <= x"c5ff4204";
		wait for Clk_period;
		Addr <=  "0010011101010";
		Trees_din <= x"00e41445";
		wait for Clk_period;
		Addr <=  "0010011101011";
		Trees_din <= x"00331445";
		wait for Clk_period;
		Addr <=  "0010011101100";
		Trees_din <= x"84fff92c";
		wait for Clk_period;
		Addr <=  "0010011101101";
		Trees_din <= x"0a00bc1c";
		wait for Clk_period;
		Addr <=  "0010011101110";
		Trees_din <= x"ccff0a0c";
		wait for Clk_period;
		Addr <=  "0010011101111";
		Trees_din <= x"0eff1f04";
		wait for Clk_period;
		Addr <=  "0010011110000";
		Trees_din <= x"ffa51445";
		wait for Clk_period;
		Addr <=  "0010011110001";
		Trees_din <= x"55004604";
		wait for Clk_period;
		Addr <=  "0010011110010";
		Trees_din <= x"00181445";
		wait for Clk_period;
		Addr <=  "0010011110011";
		Trees_din <= x"00c11445";
		wait for Clk_period;
		Addr <=  "0010011110100";
		Trees_din <= x"22019f08";
		wait for Clk_period;
		Addr <=  "0010011110101";
		Trees_din <= x"48fe8a04";
		wait for Clk_period;
		Addr <=  "0010011110110";
		Trees_din <= x"002a1445";
		wait for Clk_period;
		Addr <=  "0010011110111";
		Trees_din <= x"ff691445";
		wait for Clk_period;
		Addr <=  "0010011111000";
		Trees_din <= x"2bff8504";
		wait for Clk_period;
		Addr <=  "0010011111001";
		Trees_din <= x"00a71445";
		wait for Clk_period;
		Addr <=  "0010011111010";
		Trees_din <= x"ff9b1445";
		wait for Clk_period;
		Addr <=  "0010011111011";
		Trees_din <= x"25002c04";
		wait for Clk_period;
		Addr <=  "0010011111100";
		Trees_din <= x"ff991445";
		wait for Clk_period;
		Addr <=  "0010011111101";
		Trees_din <= x"80ff8b04";
		wait for Clk_period;
		Addr <=  "0010011111110";
		Trees_din <= x"ffbe1445";
		wait for Clk_period;
		Addr <=  "0010011111111";
		Trees_din <= x"b1fef804";
		wait for Clk_period;
		Addr <=  "0010100000000";
		Trees_din <= x"00ce1445";
		wait for Clk_period;
		Addr <=  "0010100000001";
		Trees_din <= x"000c1445";
		wait for Clk_period;
		Addr <=  "0010100000010";
		Trees_din <= x"88fff008";
		wait for Clk_period;
		Addr <=  "0010100000011";
		Trees_din <= x"dc00a004";
		wait for Clk_period;
		Addr <=  "0010100000100";
		Trees_din <= x"ff761445";
		wait for Clk_period;
		Addr <=  "0010100000101";
		Trees_din <= x"00371445";
		wait for Clk_period;
		Addr <=  "0010100000110";
		Trees_din <= x"2bff2008";
		wait for Clk_period;
		Addr <=  "0010100000111";
		Trees_din <= x"71ff3d04";
		wait for Clk_period;
		Addr <=  "0010100001000";
		Trees_din <= x"00d51445";
		wait for Clk_period;
		Addr <=  "0010100001001";
		Trees_din <= x"fffd1445";
		wait for Clk_period;
		Addr <=  "0010100001010";
		Trees_din <= x"9cffe208";
		wait for Clk_period;
		Addr <=  "0010100001011";
		Trees_din <= x"fb006704";
		wait for Clk_period;
		Addr <=  "0010100001100";
		Trees_din <= x"ffa21445";
		wait for Clk_period;
		Addr <=  "0010100001101";
		Trees_din <= x"00981445";
		wait for Clk_period;
		Addr <=  "0010100001110";
		Trees_din <= x"cbffa904";
		wait for Clk_period;
		Addr <=  "0010100001111";
		Trees_din <= x"ffd51445";
		wait for Clk_period;
		Addr <=  "0010100010000";
		Trees_din <= x"00b31445";
		wait for Clk_period;
		Addr <=  "0010100010001";
		Trees_din <= x"00ff4138";
		wait for Clk_period;
		Addr <=  "0010100010010";
		Trees_din <= x"e1000a1c";
		wait for Clk_period;
		Addr <=  "0010100010011";
		Trees_din <= x"dc00ed14";
		wait for Clk_period;
		Addr <=  "0010100010100";
		Trees_din <= x"8900a80c";
		wait for Clk_period;
		Addr <=  "0010100010101";
		Trees_din <= x"eeff0d04";
		wait for Clk_period;
		Addr <=  "0010100010110";
		Trees_din <= x"00251561";
		wait for Clk_period;
		Addr <=  "0010100010111";
		Trees_din <= x"f0002204";
		wait for Clk_period;
		Addr <=  "0010100011000";
		Trees_din <= x"ff691561";
		wait for Clk_period;
		Addr <=  "0010100011001";
		Trees_din <= x"ffee1561";
		wait for Clk_period;
		Addr <=  "0010100011010";
		Trees_din <= x"ebff5604";
		wait for Clk_period;
		Addr <=  "0010100011011";
		Trees_din <= x"ff9b1561";
		wait for Clk_period;
		Addr <=  "0010100011100";
		Trees_din <= x"007c1561";
		wait for Clk_period;
		Addr <=  "0010100011101";
		Trees_din <= x"e2fea504";
		wait for Clk_period;
		Addr <=  "0010100011110";
		Trees_din <= x"005f1561";
		wait for Clk_period;
		Addr <=  "0010100011111";
		Trees_din <= x"fff71561";
		wait for Clk_period;
		Addr <=  "0010100100000";
		Trees_din <= x"1f002f0c";
		wait for Clk_period;
		Addr <=  "0010100100001";
		Trees_din <= x"56ffe104";
		wait for Clk_period;
		Addr <=  "0010100100010";
		Trees_din <= x"ff891561";
		wait for Clk_period;
		Addr <=  "0010100100011";
		Trees_din <= x"e2fea504";
		wait for Clk_period;
		Addr <=  "0010100100100";
		Trees_din <= x"006a1561";
		wait for Clk_period;
		Addr <=  "0010100100101";
		Trees_din <= x"ffda1561";
		wait for Clk_period;
		Addr <=  "0010100100110";
		Trees_din <= x"9cff9204";
		wait for Clk_period;
		Addr <=  "0010100100111";
		Trees_din <= x"ffa41561";
		wait for Clk_period;
		Addr <=  "0010100101000";
		Trees_din <= x"0efe5904";
		wait for Clk_period;
		Addr <=  "0010100101001";
		Trees_din <= x"ffdc1561";
		wait for Clk_period;
		Addr <=  "0010100101010";
		Trees_din <= x"eeffda04";
		wait for Clk_period;
		Addr <=  "0010100101011";
		Trees_din <= x"00d71561";
		wait for Clk_period;
		Addr <=  "0010100101100";
		Trees_din <= x"00431561";
		wait for Clk_period;
		Addr <=  "0010100101101";
		Trees_din <= x"3bff3230";
		wait for Clk_period;
		Addr <=  "0010100101110";
		Trees_din <= x"71ff3418";
		wait for Clk_period;
		Addr <=  "0010100101111";
		Trees_din <= x"d2ff3810";
		wait for Clk_period;
		Addr <=  "0010100110000";
		Trees_din <= x"0fffaa08";
		wait for Clk_period;
		Addr <=  "0010100110001";
		Trees_din <= x"f7ff2404";
		wait for Clk_period;
		Addr <=  "0010100110010";
		Trees_din <= x"001d1561";
		wait for Clk_period;
		Addr <=  "0010100110011";
		Trees_din <= x"00941561";
		wait for Clk_period;
		Addr <=  "0010100110100";
		Trees_din <= x"4aff6304";
		wait for Clk_period;
		Addr <=  "0010100110101";
		Trees_din <= x"ff9e1561";
		wait for Clk_period;
		Addr <=  "0010100110110";
		Trees_din <= x"00661561";
		wait for Clk_period;
		Addr <=  "0010100110111";
		Trees_din <= x"e1008804";
		wait for Clk_period;
		Addr <=  "0010100111000";
		Trees_din <= x"ff871561";
		wait for Clk_period;
		Addr <=  "0010100111001";
		Trees_din <= x"002f1561";
		wait for Clk_period;
		Addr <=  "0010100111010";
		Trees_din <= x"11ff7d08";
		wait for Clk_period;
		Addr <=  "0010100111011";
		Trees_din <= x"6aff1904";
		wait for Clk_period;
		Addr <=  "0010100111100";
		Trees_din <= x"001f1561";
		wait for Clk_period;
		Addr <=  "0010100111101";
		Trees_din <= x"ff721561";
		wait for Clk_period;
		Addr <=  "0010100111110";
		Trees_din <= x"faffbc08";
		wait for Clk_period;
		Addr <=  "0010100111111";
		Trees_din <= x"46fece04";
		wait for Clk_period;
		Addr <=  "0010101000000";
		Trees_din <= x"005f1561";
		wait for Clk_period;
		Addr <=  "0010101000001";
		Trees_din <= x"ff9f1561";
		wait for Clk_period;
		Addr <=  "0010101000010";
		Trees_din <= x"f3feab04";
		wait for Clk_period;
		Addr <=  "0010101000011";
		Trees_din <= x"ffe81561";
		wait for Clk_period;
		Addr <=  "0010101000100";
		Trees_din <= x"009f1561";
		wait for Clk_period;
		Addr <=  "0010101000101";
		Trees_din <= x"a0fe8408";
		wait for Clk_period;
		Addr <=  "0010101000110";
		Trees_din <= x"65fe9d04";
		wait for Clk_period;
		Addr <=  "0010101000111";
		Trees_din <= x"00261561";
		wait for Clk_period;
		Addr <=  "0010101001000";
		Trees_din <= x"ff6d1561";
		wait for Clk_period;
		Addr <=  "0010101001001";
		Trees_din <= x"07005910";
		wait for Clk_period;
		Addr <=  "0010101001010";
		Trees_din <= x"53ff6a08";
		wait for Clk_period;
		Addr <=  "0010101001011";
		Trees_din <= x"53ff5a04";
		wait for Clk_period;
		Addr <=  "0010101001100";
		Trees_din <= x"ffbe1561";
		wait for Clk_period;
		Addr <=  "0010101001101";
		Trees_din <= x"00b61561";
		wait for Clk_period;
		Addr <=  "0010101001110";
		Trees_din <= x"67fe9d04";
		wait for Clk_period;
		Addr <=  "0010101001111";
		Trees_din <= x"00271561";
		wait for Clk_period;
		Addr <=  "0010101010000";
		Trees_din <= x"ff6d1561";
		wait for Clk_period;
		Addr <=  "0010101010001";
		Trees_din <= x"c5ff2808";
		wait for Clk_period;
		Addr <=  "0010101010010";
		Trees_din <= x"31fff104";
		wait for Clk_period;
		Addr <=  "0010101010011";
		Trees_din <= x"009a1561";
		wait for Clk_period;
		Addr <=  "0010101010100";
		Trees_din <= x"fff51561";
		wait for Clk_period;
		Addr <=  "0010101010101";
		Trees_din <= x"f800e004";
		wait for Clk_period;
		Addr <=  "0010101010110";
		Trees_din <= x"ffcc1561";
		wait for Clk_period;
		Addr <=  "0010101010111";
		Trees_din <= x"008f1561";
		wait for Clk_period;
		Addr <=  "0010101011000";
		Trees_din <= x"73ffd340";
		wait for Clk_period;
		Addr <=  "0010101011001";
		Trees_din <= x"82fec51c";
		wait for Clk_period;
		Addr <=  "0010101011010";
		Trees_din <= x"c5ff3110";
		wait for Clk_period;
		Addr <=  "0010101011011";
		Trees_din <= x"49000a0c";
		wait for Clk_period;
		Addr <=  "0010101011100";
		Trees_din <= x"71ff3108";
		wait for Clk_period;
		Addr <=  "0010101011101";
		Trees_din <= x"c5ff1f04";
		wait for Clk_period;
		Addr <=  "0010101011110";
		Trees_din <= x"00241695";
		wait for Clk_period;
		Addr <=  "0010101011111";
		Trees_din <= x"00d51695";
		wait for Clk_period;
		Addr <=  "0010101100000";
		Trees_din <= x"ffde1695";
		wait for Clk_period;
		Addr <=  "0010101100001";
		Trees_din <= x"ffa31695";
		wait for Clk_period;
		Addr <=  "0010101100010";
		Trees_din <= x"9dffbf04";
		wait for Clk_period;
		Addr <=  "0010101100011";
		Trees_din <= x"ff861695";
		wait for Clk_period;
		Addr <=  "0010101100100";
		Trees_din <= x"89002104";
		wait for Clk_period;
		Addr <=  "0010101100101";
		Trees_din <= x"ffcb1695";
		wait for Clk_period;
		Addr <=  "0010101100110";
		Trees_din <= x"005c1695";
		wait for Clk_period;
		Addr <=  "0010101100111";
		Trees_din <= x"8dfea408";
		wait for Clk_period;
		Addr <=  "0010101101000";
		Trees_din <= x"89017604";
		wait for Clk_period;
		Addr <=  "0010101101001";
		Trees_din <= x"ff6c1695";
		wait for Clk_period;
		Addr <=  "0010101101010";
		Trees_din <= x"00281695";
		wait for Clk_period;
		Addr <=  "0010101101011";
		Trees_din <= x"89002810";
		wait for Clk_period;
		Addr <=  "0010101101100";
		Trees_din <= x"51001408";
		wait for Clk_period;
		Addr <=  "0010101101101";
		Trees_din <= x"15003104";
		wait for Clk_period;
		Addr <=  "0010101101110";
		Trees_din <= x"ff6e1695";
		wait for Clk_period;
		Addr <=  "0010101101111";
		Trees_din <= x"00231695";
		wait for Clk_period;
		Addr <=  "0010101110000";
		Trees_din <= x"d7005604";
		wait for Clk_period;
		Addr <=  "0010101110001";
		Trees_din <= x"ff961695";
		wait for Clk_period;
		Addr <=  "0010101110010";
		Trees_din <= x"00571695";
		wait for Clk_period;
		Addr <=  "0010101110011";
		Trees_din <= x"6d000f04";
		wait for Clk_period;
		Addr <=  "0010101110100";
		Trees_din <= x"ff9f1695";
		wait for Clk_period;
		Addr <=  "0010101110101";
		Trees_din <= x"f2023104";
		wait for Clk_period;
		Addr <=  "0010101110110";
		Trees_din <= x"ffee1695";
		wait for Clk_period;
		Addr <=  "0010101110111";
		Trees_din <= x"009f1695";
		wait for Clk_period;
		Addr <=  "0010101111000";
		Trees_din <= x"39ffc43c";
		wait for Clk_period;
		Addr <=  "0010101111001";
		Trees_din <= x"30ffbe1c";
		wait for Clk_period;
		Addr <=  "0010101111010";
		Trees_din <= x"f3ff190c";
		wait for Clk_period;
		Addr <=  "0010101111011";
		Trees_din <= x"11005e08";
		wait for Clk_period;
		Addr <=  "0010101111100";
		Trees_din <= x"c2001504";
		wait for Clk_period;
		Addr <=  "0010101111101";
		Trees_din <= x"ff741695";
		wait for Clk_period;
		Addr <=  "0010101111110";
		Trees_din <= x"fff11695";
		wait for Clk_period;
		Addr <=  "0010101111111";
		Trees_din <= x"003a1695";
		wait for Clk_period;
		Addr <=  "0010110000000";
		Trees_din <= x"1effba08";
		wait for Clk_period;
		Addr <=  "0010110000001";
		Trees_din <= x"70fe5d04";
		wait for Clk_period;
		Addr <=  "0010110000010";
		Trees_din <= x"003c1695";
		wait for Clk_period;
		Addr <=  "0010110000011";
		Trees_din <= x"ff8b1695";
		wait for Clk_period;
		Addr <=  "0010110000100";
		Trees_din <= x"9cff8004";
		wait for Clk_period;
		Addr <=  "0010110000101";
		Trees_din <= x"ffe11695";
		wait for Clk_period;
		Addr <=  "0010110000110";
		Trees_din <= x"00a71695";
		wait for Clk_period;
		Addr <=  "0010110000111";
		Trees_din <= x"a3ffa510";
		wait for Clk_period;
		Addr <=  "0010110001000";
		Trees_din <= x"cf004208";
		wait for Clk_period;
		Addr <=  "0010110001001";
		Trees_din <= x"88ffe804";
		wait for Clk_period;
		Addr <=  "0010110001010";
		Trees_din <= x"ffbb1695";
		wait for Clk_period;
		Addr <=  "0010110001011";
		Trees_din <= x"006b1695";
		wait for Clk_period;
		Addr <=  "0010110001100";
		Trees_din <= x"1dfe8604";
		wait for Clk_period;
		Addr <=  "0010110001101";
		Trees_din <= x"002a1695";
		wait for Clk_period;
		Addr <=  "0010110001110";
		Trees_din <= x"ff821695";
		wait for Clk_period;
		Addr <=  "0010110001111";
		Trees_din <= x"71ff4708";
		wait for Clk_period;
		Addr <=  "0010110010000";
		Trees_din <= x"2cff3604";
		wait for Clk_period;
		Addr <=  "0010110010001";
		Trees_din <= x"ffe21695";
		wait for Clk_period;
		Addr <=  "0010110010010";
		Trees_din <= x"009c1695";
		wait for Clk_period;
		Addr <=  "0010110010011";
		Trees_din <= x"52ff0304";
		wait for Clk_period;
		Addr <=  "0010110010100";
		Trees_din <= x"004d1695";
		wait for Clk_period;
		Addr <=  "0010110010101";
		Trees_din <= x"ff9e1695";
		wait for Clk_period;
		Addr <=  "0010110010110";
		Trees_din <= x"c3001618";
		wait for Clk_period;
		Addr <=  "0010110010111";
		Trees_din <= x"2700090c";
		wait for Clk_period;
		Addr <=  "0010110011000";
		Trees_din <= x"f3ffb608";
		wait for Clk_period;
		Addr <=  "0010110011001";
		Trees_din <= x"7efdf204";
		wait for Clk_period;
		Addr <=  "0010110011010";
		Trees_din <= x"004f1695";
		wait for Clk_period;
		Addr <=  "0010110011011";
		Trees_din <= x"ff7e1695";
		wait for Clk_period;
		Addr <=  "0010110011100";
		Trees_din <= x"00831695";
		wait for Clk_period;
		Addr <=  "0010110011101";
		Trees_din <= x"80ff6404";
		wait for Clk_period;
		Addr <=  "0010110011110";
		Trees_din <= x"ffaa1695";
		wait for Clk_period;
		Addr <=  "0010110011111";
		Trees_din <= x"93ffc504";
		wait for Clk_period;
		Addr <=  "0010110100000";
		Trees_din <= x"00901695";
		wait for Clk_period;
		Addr <=  "0010110100001";
		Trees_din <= x"ffde1695";
		wait for Clk_period;
		Addr <=  "0010110100010";
		Trees_din <= x"3bffdd04";
		wait for Clk_period;
		Addr <=  "0010110100011";
		Trees_din <= x"ff721695";
		wait for Clk_period;
		Addr <=  "0010110100100";
		Trees_din <= x"fff91695";
		wait for Clk_period;
		Addr <=  "0010110100101";
		Trees_din <= x"9cff9454";
		wait for Clk_period;
		Addr <=  "0010110100110";
		Trees_din <= x"0a004a20";
		wait for Clk_period;
		Addr <=  "0010110100111";
		Trees_din <= x"2e006b18";
		wait for Clk_period;
		Addr <=  "0010110101000";
		Trees_din <= x"18013b0c";
		wait for Clk_period;
		Addr <=  "0010110101001";
		Trees_din <= x"ab015008";
		wait for Clk_period;
		Addr <=  "0010110101010";
		Trees_din <= x"43fed904";
		wait for Clk_period;
		Addr <=  "0010110101011";
		Trees_din <= x"ffdf17f1";
		wait for Clk_period;
		Addr <=  "0010110101100";
		Trees_din <= x"ff7017f1";
		wait for Clk_period;
		Addr <=  "0010110101101";
		Trees_din <= x"003817f1";
		wait for Clk_period;
		Addr <=  "0010110101110";
		Trees_din <= x"baffb008";
		wait for Clk_period;
		Addr <=  "0010110101111";
		Trees_din <= x"f1ff6704";
		wait for Clk_period;
		Addr <=  "0010110110000";
		Trees_din <= x"009f17f1";
		wait for Clk_period;
		Addr <=  "0010110110001";
		Trees_din <= x"ffeb17f1";
		wait for Clk_period;
		Addr <=  "0010110110010";
		Trees_din <= x"ff9d17f1";
		wait for Clk_period;
		Addr <=  "0010110110011";
		Trees_din <= x"62fedf04";
		wait for Clk_period;
		Addr <=  "0010110110100";
		Trees_din <= x"009217f1";
		wait for Clk_period;
		Addr <=  "0010110110101";
		Trees_din <= x"ffe817f1";
		wait for Clk_period;
		Addr <=  "0010110110110";
		Trees_din <= x"8e00411c";
		wait for Clk_period;
		Addr <=  "0010110110111";
		Trees_din <= x"bcfeb110";
		wait for Clk_period;
		Addr <=  "0010110111000";
		Trees_din <= x"f0ff4008";
		wait for Clk_period;
		Addr <=  "0010110111001";
		Trees_din <= x"47002504";
		wait for Clk_period;
		Addr <=  "0010110111010";
		Trees_din <= x"ffdd17f1";
		wait for Clk_period;
		Addr <=  "0010110111011";
		Trees_din <= x"007e17f1";
		wait for Clk_period;
		Addr <=  "0010110111100";
		Trees_din <= x"a6ff1504";
		wait for Clk_period;
		Addr <=  "0010110111101";
		Trees_din <= x"002017f1";
		wait for Clk_period;
		Addr <=  "0010110111110";
		Trees_din <= x"ff9e17f1";
		wait for Clk_period;
		Addr <=  "0010110111111";
		Trees_din <= x"ddffb308";
		wait for Clk_period;
		Addr <=  "0010111000000";
		Trees_din <= x"77002404";
		wait for Clk_period;
		Addr <=  "0010111000001";
		Trees_din <= x"ff7317f1";
		wait for Clk_period;
		Addr <=  "0010111000010";
		Trees_din <= x"000317f1";
		wait for Clk_period;
		Addr <=  "0010111000011";
		Trees_din <= x"006c17f1";
		wait for Clk_period;
		Addr <=  "0010111000100";
		Trees_din <= x"a8ffd910";
		wait for Clk_period;
		Addr <=  "0010111000101";
		Trees_din <= x"2cffa708";
		wait for Clk_period;
		Addr <=  "0010111000110";
		Trees_din <= x"7fffe104";
		wait for Clk_period;
		Addr <=  "0010111000111";
		Trees_din <= x"ffa017f1";
		wait for Clk_period;
		Addr <=  "0010111001000";
		Trees_din <= x"006517f1";
		wait for Clk_period;
		Addr <=  "0010111001001";
		Trees_din <= x"15ff7504";
		wait for Clk_period;
		Addr <=  "0010111001010";
		Trees_din <= x"00a117f1";
		wait for Clk_period;
		Addr <=  "0010111001011";
		Trees_din <= x"001b17f1";
		wait for Clk_period;
		Addr <=  "0010111001100";
		Trees_din <= x"e7ff7304";
		wait for Clk_period;
		Addr <=  "0010111001101";
		Trees_din <= x"ffe217f1";
		wait for Clk_period;
		Addr <=  "0010111001110";
		Trees_din <= x"ff9217f1";
		wait for Clk_period;
		Addr <=  "0010111001111";
		Trees_din <= x"73ffbd24";
		wait for Clk_period;
		Addr <=  "0010111010000";
		Trees_din <= x"82ff0b14";
		wait for Clk_period;
		Addr <=  "0010111010001";
		Trees_din <= x"56ff6010";
		wait for Clk_period;
		Addr <=  "0010111010010";
		Trees_din <= x"5dffaf08";
		wait for Clk_period;
		Addr <=  "0010111010011";
		Trees_din <= x"78ff5f04";
		wait for Clk_period;
		Addr <=  "0010111010100";
		Trees_din <= x"001617f1";
		wait for Clk_period;
		Addr <=  "0010111010101";
		Trees_din <= x"00ab17f1";
		wait for Clk_period;
		Addr <=  "0010111010110";
		Trees_din <= x"d2feee04";
		wait for Clk_period;
		Addr <=  "0010111010111";
		Trees_din <= x"ffb017f1";
		wait for Clk_period;
		Addr <=  "0010111011000";
		Trees_din <= x"001217f1";
		wait for Clk_period;
		Addr <=  "0010111011001";
		Trees_din <= x"ffa117f1";
		wait for Clk_period;
		Addr <=  "0010111011010";
		Trees_din <= x"d6008b04";
		wait for Clk_period;
		Addr <=  "0010111011011";
		Trees_din <= x"ff7217f1";
		wait for Clk_period;
		Addr <=  "0010111011100";
		Trees_din <= x"54006c04";
		wait for Clk_period;
		Addr <=  "0010111011101";
		Trees_din <= x"ffa817f1";
		wait for Clk_period;
		Addr <=  "0010111011110";
		Trees_din <= x"dfff8704";
		wait for Clk_period;
		Addr <=  "0010111011111";
		Trees_din <= x"001117f1";
		wait for Clk_period;
		Addr <=  "0010111100000";
		Trees_din <= x"006317f1";
		wait for Clk_period;
		Addr <=  "0010111100001";
		Trees_din <= x"28ff2918";
		wait for Clk_period;
		Addr <=  "0010111100010";
		Trees_din <= x"10ff0e08";
		wait for Clk_period;
		Addr <=  "0010111100011";
		Trees_din <= x"78ffca04";
		wait for Clk_period;
		Addr <=  "0010111100100";
		Trees_din <= x"ffff17f1";
		wait for Clk_period;
		Addr <=  "0010111100101";
		Trees_din <= x"00a217f1";
		wait for Clk_period;
		Addr <=  "0010111100110";
		Trees_din <= x"01fe3a08";
		wait for Clk_period;
		Addr <=  "0010111100111";
		Trees_din <= x"00ffde04";
		wait for Clk_period;
		Addr <=  "0010111101000";
		Trees_din <= x"ffd517f1";
		wait for Clk_period;
		Addr <=  "0010111101001";
		Trees_din <= x"007017f1";
		wait for Clk_period;
		Addr <=  "0010111101010";
		Trees_din <= x"11000804";
		wait for Clk_period;
		Addr <=  "0010111101011";
		Trees_din <= x"ff7817f1";
		wait for Clk_period;
		Addr <=  "0010111101100";
		Trees_din <= x"001117f1";
		wait for Clk_period;
		Addr <=  "0010111101101";
		Trees_din <= x"89ff7d10";
		wait for Clk_period;
		Addr <=  "0010111101110";
		Trees_din <= x"17ffec08";
		wait for Clk_period;
		Addr <=  "0010111101111";
		Trees_din <= x"a6ffb004";
		wait for Clk_period;
		Addr <=  "0010111110000";
		Trees_din <= x"ffe917f1";
		wait for Clk_period;
		Addr <=  "0010111110001";
		Trees_din <= x"006517f1";
		wait for Clk_period;
		Addr <=  "0010111110010";
		Trees_din <= x"d6006504";
		wait for Clk_period;
		Addr <=  "0010111110011";
		Trees_din <= x"00ef17f1";
		wait for Clk_period;
		Addr <=  "0010111110100";
		Trees_din <= x"004217f1";
		wait for Clk_period;
		Addr <=  "0010111110101";
		Trees_din <= x"e8ff6608";
		wait for Clk_period;
		Addr <=  "0010111110110";
		Trees_din <= x"e1ffd004";
		wait for Clk_period;
		Addr <=  "0010111110111";
		Trees_din <= x"ffe517f1";
		wait for Clk_period;
		Addr <=  "0010111111000";
		Trees_din <= x"008617f1";
		wait for Clk_period;
		Addr <=  "0010111111001";
		Trees_din <= x"baffc804";
		wait for Clk_period;
		Addr <=  "0010111111010";
		Trees_din <= x"ff8c17f1";
		wait for Clk_period;
		Addr <=  "0010111111011";
		Trees_din <= x"003e17f1";
		wait for Clk_period;
		Addr <=  "0010111111100";
		Trees_din <= x"8dfe9040";
		wait for Clk_period;
		Addr <=  "0010111111101";
		Trees_din <= x"73ffd514";
		wait for Clk_period;
		Addr <=  "0010111111110";
		Trees_din <= x"3afeb610";
		wait for Clk_period;
		Addr <=  "0010111111111";
		Trees_din <= x"f3ff0904";
		wait for Clk_period;
		Addr <=  "0011000000000";
		Trees_din <= x"ff8e193d";
		wait for Clk_period;
		Addr <=  "0011000000001";
		Trees_din <= x"cbffbc04";
		wait for Clk_period;
		Addr <=  "0011000000010";
		Trees_din <= x"ffc6193d";
		wait for Clk_period;
		Addr <=  "0011000000011";
		Trees_din <= x"9bff0704";
		wait for Clk_period;
		Addr <=  "0011000000100";
		Trees_din <= x"0078193d";
		wait for Clk_period;
		Addr <=  "0011000000101";
		Trees_din <= x"0009193d";
		wait for Clk_period;
		Addr <=  "0011000000110";
		Trees_din <= x"ff72193d";
		wait for Clk_period;
		Addr <=  "0011000000111";
		Trees_din <= x"68fe9618";
		wait for Clk_period;
		Addr <=  "0011000001000";
		Trees_din <= x"f7ff4608";
		wait for Clk_period;
		Addr <=  "0011000001001";
		Trees_din <= x"69fe8904";
		wait for Clk_period;
		Addr <=  "0011000001010";
		Trees_din <= x"0040193d";
		wait for Clk_period;
		Addr <=  "0011000001011";
		Trees_din <= x"ff91193d";
		wait for Clk_period;
		Addr <=  "0011000001100";
		Trees_din <= x"27fff808";
		wait for Clk_period;
		Addr <=  "0011000001101";
		Trees_din <= x"8dfe6104";
		wait for Clk_period;
		Addr <=  "0011000001110";
		Trees_din <= x"ffb4193d";
		wait for Clk_period;
		Addr <=  "0011000001111";
		Trees_din <= x"004d193d";
		wait for Clk_period;
		Addr <=  "0011000010000";
		Trees_din <= x"7dffe904";
		wait for Clk_period;
		Addr <=  "0011000010001";
		Trees_din <= x"00ac193d";
		wait for Clk_period;
		Addr <=  "0011000010010";
		Trees_din <= x"001a193d";
		wait for Clk_period;
		Addr <=  "0011000010011";
		Trees_din <= x"d4ff1804";
		wait for Clk_period;
		Addr <=  "0011000010100";
		Trees_din <= x"ff77193d";
		wait for Clk_period;
		Addr <=  "0011000010101";
		Trees_din <= x"7d003808";
		wait for Clk_period;
		Addr <=  "0011000010110";
		Trees_din <= x"72ffb404";
		wait for Clk_period;
		Addr <=  "0011000010111";
		Trees_din <= x"0041193d";
		wait for Clk_period;
		Addr <=  "0011000011000";
		Trees_din <= x"ff96193d";
		wait for Clk_period;
		Addr <=  "0011000011001";
		Trees_din <= x"d000be04";
		wait for Clk_period;
		Addr <=  "0011000011010";
		Trees_din <= x"ffd4193d";
		wait for Clk_period;
		Addr <=  "0011000011011";
		Trees_din <= x"006d193d";
		wait for Clk_period;
		Addr <=  "0011000011100";
		Trees_din <= x"1afec138";
		wait for Clk_period;
		Addr <=  "0011000011101";
		Trees_din <= x"66ffac18";
		wait for Clk_period;
		Addr <=  "0011000011110";
		Trees_din <= x"baff9710";
		wait for Clk_period;
		Addr <=  "0011000011111";
		Trees_din <= x"79ff5308";
		wait for Clk_period;
		Addr <=  "0011000100000";
		Trees_din <= x"32fead04";
		wait for Clk_period;
		Addr <=  "0011000100001";
		Trees_din <= x"ffd3193d";
		wait for Clk_period;
		Addr <=  "0011000100010";
		Trees_din <= x"0075193d";
		wait for Clk_period;
		Addr <=  "0011000100011";
		Trees_din <= x"6d003104";
		wait for Clk_period;
		Addr <=  "0011000100100";
		Trees_din <= x"ffa5193d";
		wait for Clk_period;
		Addr <=  "0011000100101";
		Trees_din <= x"ffec193d";
		wait for Clk_period;
		Addr <=  "0011000100110";
		Trees_din <= x"11ffec04";
		wait for Clk_period;
		Addr <=  "0011000100111";
		Trees_din <= x"ff81193d";
		wait for Clk_period;
		Addr <=  "0011000101000";
		Trees_din <= x"fffb193d";
		wait for Clk_period;
		Addr <=  "0011000101001";
		Trees_din <= x"cbffe210";
		wait for Clk_period;
		Addr <=  "0011000101010";
		Trees_din <= x"f7003a08";
		wait for Clk_period;
		Addr <=  "0011000101011";
		Trees_din <= x"8ffe5904";
		wait for Clk_period;
		Addr <=  "0011000101100";
		Trees_din <= x"ffd3193d";
		wait for Clk_period;
		Addr <=  "0011000101101";
		Trees_din <= x"0084193d";
		wait for Clk_period;
		Addr <=  "0011000101110";
		Trees_din <= x"d1ff1b04";
		wait for Clk_period;
		Addr <=  "0011000101111";
		Trees_din <= x"0031193d";
		wait for Clk_period;
		Addr <=  "0011000110000";
		Trees_din <= x"ff9c193d";
		wait for Clk_period;
		Addr <=  "0011000110001";
		Trees_din <= x"90fffe08";
		wait for Clk_period;
		Addr <=  "0011000110010";
		Trees_din <= x"c4fe6404";
		wait for Clk_period;
		Addr <=  "0011000110011";
		Trees_din <= x"0034193d";
		wait for Clk_period;
		Addr <=  "0011000110100";
		Trees_din <= x"ff82193d";
		wait for Clk_period;
		Addr <=  "0011000110101";
		Trees_din <= x"1afe2404";
		wait for Clk_period;
		Addr <=  "0011000110110";
		Trees_din <= x"007b193d";
		wait for Clk_period;
		Addr <=  "0011000110111";
		Trees_din <= x"ffeb193d";
		wait for Clk_period;
		Addr <=  "0011000111000";
		Trees_din <= x"93ffd018";
		wait for Clk_period;
		Addr <=  "0011000111001";
		Trees_din <= x"8900c510";
		wait for Clk_period;
		Addr <=  "0011000111010";
		Trees_din <= x"08004f08";
		wait for Clk_period;
		Addr <=  "0011000111011";
		Trees_din <= x"9bffee04";
		wait for Clk_period;
		Addr <=  "0011000111100";
		Trees_din <= x"ff6f193d";
		wait for Clk_period;
		Addr <=  "0011000111101";
		Trees_din <= x"fffc193d";
		wait for Clk_period;
		Addr <=  "0011000111110";
		Trees_din <= x"a9ff7404";
		wait for Clk_period;
		Addr <=  "0011000111111";
		Trees_din <= x"0029193d";
		wait for Clk_period;
		Addr <=  "0011001000000";
		Trees_din <= x"ff9a193d";
		wait for Clk_period;
		Addr <=  "0011001000001";
		Trees_din <= x"a5fed704";
		wait for Clk_period;
		Addr <=  "0011001000010";
		Trees_din <= x"0086193d";
		wait for Clk_period;
		Addr <=  "0011001000011";
		Trees_din <= x"0019193d";
		wait for Clk_period;
		Addr <=  "0011001000100";
		Trees_din <= x"02fe5e08";
		wait for Clk_period;
		Addr <=  "0011001000101";
		Trees_din <= x"c7fee604";
		wait for Clk_period;
		Addr <=  "0011001000110";
		Trees_din <= x"00bb193d";
		wait for Clk_period;
		Addr <=  "0011001000111";
		Trees_din <= x"0020193d";
		wait for Clk_period;
		Addr <=  "0011001001000";
		Trees_din <= x"a6ff8708";
		wait for Clk_period;
		Addr <=  "0011001001001";
		Trees_din <= x"c6ff1304";
		wait for Clk_period;
		Addr <=  "0011001001010";
		Trees_din <= x"0021193d";
		wait for Clk_period;
		Addr <=  "0011001001011";
		Trees_din <= x"ff85193d";
		wait for Clk_period;
		Addr <=  "0011001001100";
		Trees_din <= x"d7009c04";
		wait for Clk_period;
		Addr <=  "0011001001101";
		Trees_din <= x"ffe9193d";
		wait for Clk_period;
		Addr <=  "0011001001110";
		Trees_din <= x"009d193d";
		wait for Clk_period;
		Addr <=  "0011001001111";
		Trees_din <= x"2fff7e50";
		wait for Clk_period;
		Addr <=  "0011001010000";
		Trees_din <= x"e6ff9f2c";
		wait for Clk_period;
		Addr <=  "0011001010001";
		Trees_din <= x"5a003718";
		wait for Clk_period;
		Addr <=  "0011001010010";
		Trees_din <= x"bbff5a0c";
		wait for Clk_period;
		Addr <=  "0011001010011";
		Trees_din <= x"bbfee008";
		wait for Clk_period;
		Addr <=  "0011001010100";
		Trees_din <= x"ebff0204";
		wait for Clk_period;
		Addr <=  "0011001010101";
		Trees_din <= x"ffe61a99";
		wait for Clk_period;
		Addr <=  "0011001010110";
		Trees_din <= x"00641a99";
		wait for Clk_period;
		Addr <=  "0011001010111";
		Trees_din <= x"ff991a99";
		wait for Clk_period;
		Addr <=  "0011001011000";
		Trees_din <= x"e6ff4504";
		wait for Clk_period;
		Addr <=  "0011001011001";
		Trees_din <= x"ffe71a99";
		wait for Clk_period;
		Addr <=  "0011001011010";
		Trees_din <= x"6fff5204";
		wait for Clk_period;
		Addr <=  "0011001011011";
		Trees_din <= x"009e1a99";
		wait for Clk_period;
		Addr <=  "0011001011100";
		Trees_din <= x"00101a99";
		wait for Clk_period;
		Addr <=  "0011001011101";
		Trees_din <= x"bdffbc10";
		wait for Clk_period;
		Addr <=  "0011001011110";
		Trees_din <= x"efff6908";
		wait for Clk_period;
		Addr <=  "0011001011111";
		Trees_din <= x"0a003a04";
		wait for Clk_period;
		Addr <=  "0011001100000";
		Trees_din <= x"ffab1a99";
		wait for Clk_period;
		Addr <=  "0011001100001";
		Trees_din <= x"00601a99";
		wait for Clk_period;
		Addr <=  "0011001100010";
		Trees_din <= x"a1ff9b04";
		wait for Clk_period;
		Addr <=  "0011001100011";
		Trees_din <= x"ff8d1a99";
		wait for Clk_period;
		Addr <=  "0011001100100";
		Trees_din <= x"00211a99";
		wait for Clk_period;
		Addr <=  "0011001100101";
		Trees_din <= x"ff761a99";
		wait for Clk_period;
		Addr <=  "0011001100110";
		Trees_din <= x"ccff0308";
		wait for Clk_period;
		Addr <=  "0011001100111";
		Trees_din <= x"3afef404";
		wait for Clk_period;
		Addr <=  "0011001101000";
		Trees_din <= x"006f1a99";
		wait for Clk_period;
		Addr <=  "0011001101001";
		Trees_din <= x"ffe31a99";
		wait for Clk_period;
		Addr <=  "0011001101010";
		Trees_din <= x"fb00080c";
		wait for Clk_period;
		Addr <=  "0011001101011";
		Trees_din <= x"0a014908";
		wait for Clk_period;
		Addr <=  "0011001101100";
		Trees_din <= x"5100e704";
		wait for Clk_period;
		Addr <=  "0011001101101";
		Trees_din <= x"ff6c1a99";
		wait for Clk_period;
		Addr <=  "0011001101110";
		Trees_din <= x"ffea1a99";
		wait for Clk_period;
		Addr <=  "0011001101111";
		Trees_din <= x"002e1a99";
		wait for Clk_period;
		Addr <=  "0011001110000";
		Trees_din <= x"bfff2408";
		wait for Clk_period;
		Addr <=  "0011001110001";
		Trees_din <= x"76001204";
		wait for Clk_period;
		Addr <=  "0011001110010";
		Trees_din <= x"ffee1a99";
		wait for Clk_period;
		Addr <=  "0011001110011";
		Trees_din <= x"00831a99";
		wait for Clk_period;
		Addr <=  "0011001110100";
		Trees_din <= x"d3feb504";
		wait for Clk_period;
		Addr <=  "0011001110101";
		Trees_din <= x"fffe1a99";
		wait for Clk_period;
		Addr <=  "0011001110110";
		Trees_din <= x"ff901a99";
		wait for Clk_period;
		Addr <=  "0011001110111";
		Trees_din <= x"67ff6638";
		wait for Clk_period;
		Addr <=  "0011001111000";
		Trees_din <= x"aaff7318";
		wait for Clk_period;
		Addr <=  "0011001111001";
		Trees_din <= x"0800950c";
		wait for Clk_period;
		Addr <=  "0011001111010";
		Trees_din <= x"a0ffb508";
		wait for Clk_period;
		Addr <=  "0011001111011";
		Trees_din <= x"fe005d04";
		wait for Clk_period;
		Addr <=  "0011001111100";
		Trees_din <= x"ff771a99";
		wait for Clk_period;
		Addr <=  "0011001111101";
		Trees_din <= x"00111a99";
		wait for Clk_period;
		Addr <=  "0011001111110";
		Trees_din <= x"00501a99";
		wait for Clk_period;
		Addr <=  "0011001111111";
		Trees_din <= x"8c009908";
		wait for Clk_period;
		Addr <=  "0011010000000";
		Trees_din <= x"9cff4904";
		wait for Clk_period;
		Addr <=  "0011010000001";
		Trees_din <= x"ffca1a99";
		wait for Clk_period;
		Addr <=  "0011010000010";
		Trees_din <= x"00741a99";
		wait for Clk_period;
		Addr <=  "0011010000011";
		Trees_din <= x"ff9f1a99";
		wait for Clk_period;
		Addr <=  "0011010000100";
		Trees_din <= x"24ffc610";
		wait for Clk_period;
		Addr <=  "0011010000101";
		Trees_din <= x"68fe9408";
		wait for Clk_period;
		Addr <=  "0011010000110";
		Trees_din <= x"2affb004";
		wait for Clk_period;
		Addr <=  "0011010000111";
		Trees_din <= x"00051a99";
		wait for Clk_period;
		Addr <=  "0011010001000";
		Trees_din <= x"00b41a99";
		wait for Clk_period;
		Addr <=  "0011010001001";
		Trees_din <= x"3bff3204";
		wait for Clk_period;
		Addr <=  "0011010001010";
		Trees_din <= x"00691a99";
		wait for Clk_period;
		Addr <=  "0011010001011";
		Trees_din <= x"ffdf1a99";
		wait for Clk_period;
		Addr <=  "0011010001100";
		Trees_din <= x"ddfec508";
		wait for Clk_period;
		Addr <=  "0011010001101";
		Trees_din <= x"02fe5204";
		wait for Clk_period;
		Addr <=  "0011010001110";
		Trees_din <= x"007f1a99";
		wait for Clk_period;
		Addr <=  "0011010001111";
		Trees_din <= x"001b1a99";
		wait for Clk_period;
		Addr <=  "0011010010000";
		Trees_din <= x"2f002404";
		wait for Clk_period;
		Addr <=  "0011010010001";
		Trees_din <= x"ff8e1a99";
		wait for Clk_period;
		Addr <=  "0011010010010";
		Trees_din <= x"001e1a99";
		wait for Clk_period;
		Addr <=  "0011010010011";
		Trees_din <= x"cd002418";
		wait for Clk_period;
		Addr <=  "0011010010100";
		Trees_din <= x"83ff1510";
		wait for Clk_period;
		Addr <=  "0011010010101";
		Trees_din <= x"1f000c08";
		wait for Clk_period;
		Addr <=  "0011010010110";
		Trees_din <= x"38fee404";
		wait for Clk_period;
		Addr <=  "0011010010111";
		Trees_din <= x"001a1a99";
		wait for Clk_period;
		Addr <=  "0011010011000";
		Trees_din <= x"ff901a99";
		wait for Clk_period;
		Addr <=  "0011010011001";
		Trees_din <= x"6bfed004";
		wait for Clk_period;
		Addr <=  "0011010011010";
		Trees_din <= x"ffe01a99";
		wait for Clk_period;
		Addr <=  "0011010011011";
		Trees_din <= x"00781a99";
		wait for Clk_period;
		Addr <=  "0011010011100";
		Trees_din <= x"fcfeb904";
		wait for Clk_period;
		Addr <=  "0011010011101";
		Trees_din <= x"00071a99";
		wait for Clk_period;
		Addr <=  "0011010011110";
		Trees_din <= x"ff741a99";
		wait for Clk_period;
		Addr <=  "0011010011111";
		Trees_din <= x"9dff9104";
		wait for Clk_period;
		Addr <=  "0011010100000";
		Trees_din <= x"ffb81a99";
		wait for Clk_period;
		Addr <=  "0011010100001";
		Trees_din <= x"40001308";
		wait for Clk_period;
		Addr <=  "0011010100010";
		Trees_din <= x"d3ff2504";
		wait for Clk_period;
		Addr <=  "0011010100011";
		Trees_din <= x"001e1a99";
		wait for Clk_period;
		Addr <=  "0011010100100";
		Trees_din <= x"009d1a99";
		wait for Clk_period;
		Addr <=  "0011010100101";
		Trees_din <= x"ffff1a99";
		wait for Clk_period;
		Addr <=  "0011010100110";
		Trees_din <= x"0fff3138";
		wait for Clk_period;
		Addr <=  "0011010100111";
		Trees_din <= x"1cff6a1c";
		wait for Clk_period;
		Addr <=  "0011010101000";
		Trees_din <= x"67ffae14";
		wait for Clk_period;
		Addr <=  "0011010101001";
		Trees_din <= x"19ff8a10";
		wait for Clk_period;
		Addr <=  "0011010101010";
		Trees_din <= x"e2ff7c08";
		wait for Clk_period;
		Addr <=  "0011010101011";
		Trees_din <= x"f7feb504";
		wait for Clk_period;
		Addr <=  "0011010101100";
		Trees_din <= x"ffde1b95";
		wait for Clk_period;
		Addr <=  "0011010101101";
		Trees_din <= x"00791b95";
		wait for Clk_period;
		Addr <=  "0011010101110";
		Trees_din <= x"e6ff7b04";
		wait for Clk_period;
		Addr <=  "0011010101111";
		Trees_din <= x"003d1b95";
		wait for Clk_period;
		Addr <=  "0011010110000";
		Trees_din <= x"ffae1b95";
		wait for Clk_period;
		Addr <=  "0011010110001";
		Trees_din <= x"ffc81b95";
		wait for Clk_period;
		Addr <=  "0011010110010";
		Trees_din <= x"43ffc304";
		wait for Clk_period;
		Addr <=  "0011010110011";
		Trees_din <= x"ff991b95";
		wait for Clk_period;
		Addr <=  "0011010110100";
		Trees_din <= x"00121b95";
		wait for Clk_period;
		Addr <=  "0011010110101";
		Trees_din <= x"11fff010";
		wait for Clk_period;
		Addr <=  "0011010110110";
		Trees_din <= x"60fef404";
		wait for Clk_period;
		Addr <=  "0011010110111";
		Trees_din <= x"00301b95";
		wait for Clk_period;
		Addr <=  "0011010111000";
		Trees_din <= x"0700e408";
		wait for Clk_period;
		Addr <=  "0011010111001";
		Trees_din <= x"f2011704";
		wait for Clk_period;
		Addr <=  "0011010111010";
		Trees_din <= x"ffe91b95";
		wait for Clk_period;
		Addr <=  "0011010111011";
		Trees_din <= x"ff771b95";
		wait for Clk_period;
		Addr <=  "0011010111100";
		Trees_din <= x"00391b95";
		wait for Clk_period;
		Addr <=  "0011010111101";
		Trees_din <= x"aeff3c08";
		wait for Clk_period;
		Addr <=  "0011010111110";
		Trees_din <= x"73000604";
		wait for Clk_period;
		Addr <=  "0011010111111";
		Trees_din <= x"00081b95";
		wait for Clk_period;
		Addr <=  "0011011000000";
		Trees_din <= x"00731b95";
		wait for Clk_period;
		Addr <=  "0011011000001";
		Trees_din <= x"ffd01b95";
		wait for Clk_period;
		Addr <=  "0011011000010";
		Trees_din <= x"30ffb518";
		wait for Clk_period;
		Addr <=  "0011011000011";
		Trees_din <= x"2c006810";
		wait for Clk_period;
		Addr <=  "0011011000100";
		Trees_din <= x"5cff6908";
		wait for Clk_period;
		Addr <=  "0011011000101";
		Trees_din <= x"b0fef104";
		wait for Clk_period;
		Addr <=  "0011011000110";
		Trees_din <= x"00691b95";
		wait for Clk_period;
		Addr <=  "0011011000111";
		Trees_din <= x"ffa61b95";
		wait for Clk_period;
		Addr <=  "0011011001000";
		Trees_din <= x"cd008504";
		wait for Clk_period;
		Addr <=  "0011011001001";
		Trees_din <= x"ff6e1b95";
		wait for Clk_period;
		Addr <=  "0011011001010";
		Trees_din <= x"ffee1b95";
		wait for Clk_period;
		Addr <=  "0011011001011";
		Trees_din <= x"c1feec04";
		wait for Clk_period;
		Addr <=  "0011011001100";
		Trees_din <= x"00061b95";
		wait for Clk_period;
		Addr <=  "0011011001101";
		Trees_din <= x"004d1b95";
		wait for Clk_period;
		Addr <=  "0011011001110";
		Trees_din <= x"a9ffac20";
		wait for Clk_period;
		Addr <=  "0011011001111";
		Trees_din <= x"2affdf10";
		wait for Clk_period;
		Addr <=  "0011011010000";
		Trees_din <= x"eeff5908";
		wait for Clk_period;
		Addr <=  "0011011010001";
		Trees_din <= x"d3ff4204";
		wait for Clk_period;
		Addr <=  "0011011010010";
		Trees_din <= x"ffec1b95";
		wait for Clk_period;
		Addr <=  "0011011010011";
		Trees_din <= x"00741b95";
		wait for Clk_period;
		Addr <=  "0011011010100";
		Trees_din <= x"6bfe2304";
		wait for Clk_period;
		Addr <=  "0011011010101";
		Trees_din <= x"00341b95";
		wait for Clk_period;
		Addr <=  "0011011010110";
		Trees_din <= x"ff931b95";
		wait for Clk_period;
		Addr <=  "0011011010111";
		Trees_din <= x"88ffd008";
		wait for Clk_period;
		Addr <=  "0011011011000";
		Trees_din <= x"d3fe9e04";
		wait for Clk_period;
		Addr <=  "0011011011001";
		Trees_din <= x"00131b95";
		wait for Clk_period;
		Addr <=  "0011011011010";
		Trees_din <= x"ff8b1b95";
		wait for Clk_period;
		Addr <=  "0011011011011";
		Trees_din <= x"31007e04";
		wait for Clk_period;
		Addr <=  "0011011011100";
		Trees_din <= x"005b1b95";
		wait for Clk_period;
		Addr <=  "0011011011101";
		Trees_din <= x"ffb81b95";
		wait for Clk_period;
		Addr <=  "0011011011110";
		Trees_din <= x"2e00810c";
		wait for Clk_period;
		Addr <=  "0011011011111";
		Trees_din <= x"55ff8b04";
		wait for Clk_period;
		Addr <=  "0011011100000";
		Trees_din <= x"00131b95";
		wait for Clk_period;
		Addr <=  "0011011100001";
		Trees_din <= x"ccff2404";
		wait for Clk_period;
		Addr <=  "0011011100010";
		Trees_din <= x"ffee1b95";
		wait for Clk_period;
		Addr <=  "0011011100011";
		Trees_din <= x"ff701b95";
		wait for Clk_period;
		Addr <=  "0011011100100";
		Trees_din <= x"00801b95";
		wait for Clk_period;
		Addr <=  "0011011100101";
		Trees_din <= x"00ff4128";
		wait for Clk_period;
		Addr <=  "0011011100110";
		Trees_din <= x"1f002f10";
		wait for Clk_period;
		Addr <=  "0011011100111";
		Trees_din <= x"ed007a0c";
		wait for Clk_period;
		Addr <=  "0011011101000";
		Trees_din <= x"4e000f08";
		wait for Clk_period;
		Addr <=  "0011011101001";
		Trees_din <= x"b8fed204";
		wait for Clk_period;
		Addr <=  "0011011101010";
		Trees_din <= x"ffda1c89";
		wait for Clk_period;
		Addr <=  "0011011101011";
		Trees_din <= x"ff701c89";
		wait for Clk_period;
		Addr <=  "0011011101100";
		Trees_din <= x"000d1c89";
		wait for Clk_period;
		Addr <=  "0011011101101";
		Trees_din <= x"002a1c89";
		wait for Clk_period;
		Addr <=  "0011011101110";
		Trees_din <= x"51ffef08";
		wait for Clk_period;
		Addr <=  "0011011101111";
		Trees_din <= x"4afe8c04";
		wait for Clk_period;
		Addr <=  "0011011110000";
		Trees_din <= x"001a1c89";
		wait for Clk_period;
		Addr <=  "0011011110001";
		Trees_din <= x"ff8c1c89";
		wait for Clk_period;
		Addr <=  "0011011110010";
		Trees_din <= x"5effbc04";
		wait for Clk_period;
		Addr <=  "0011011110011";
		Trees_din <= x"ffcd1c89";
		wait for Clk_period;
		Addr <=  "0011011110100";
		Trees_din <= x"2a000b08";
		wait for Clk_period;
		Addr <=  "0011011110101";
		Trees_din <= x"76ffa404";
		wait for Clk_period;
		Addr <=  "0011011110110";
		Trees_din <= x"00991c89";
		wait for Clk_period;
		Addr <=  "0011011110111";
		Trees_din <= x"00211c89";
		wait for Clk_period;
		Addr <=  "0011011111000";
		Trees_din <= x"000f1c89";
		wait for Clk_period;
		Addr <=  "0011011111001";
		Trees_din <= x"24ffe034";
		wait for Clk_period;
		Addr <=  "0011011111010";
		Trees_din <= x"4bff101c";
		wait for Clk_period;
		Addr <=  "0011011111011";
		Trees_din <= x"2fff8c10";
		wait for Clk_period;
		Addr <=  "0011011111100";
		Trees_din <= x"c7feff08";
		wait for Clk_period;
		Addr <=  "0011011111101";
		Trees_din <= x"8dfe6404";
		wait for Clk_period;
		Addr <=  "0011011111110";
		Trees_din <= x"ffc91c89";
		wait for Clk_period;
		Addr <=  "0011011111111";
		Trees_din <= x"003d1c89";
		wait for Clk_period;
		Addr <=  "0011100000000";
		Trees_din <= x"00ffd904";
		wait for Clk_period;
		Addr <=  "0011100000001";
		Trees_din <= x"ff801c89";
		wait for Clk_period;
		Addr <=  "0011100000010";
		Trees_din <= x"00241c89";
		wait for Clk_period;
		Addr <=  "0011100000011";
		Trees_din <= x"2aff8804";
		wait for Clk_period;
		Addr <=  "0011100000100";
		Trees_din <= x"ffc51c89";
		wait for Clk_period;
		Addr <=  "0011100000101";
		Trees_din <= x"87ff2b04";
		wait for Clk_period;
		Addr <=  "0011100000110";
		Trees_din <= x"00011c89";
		wait for Clk_period;
		Addr <=  "0011100000111";
		Trees_din <= x"006c1c89";
		wait for Clk_period;
		Addr <=  "0011100001000";
		Trees_din <= x"28ff9f10";
		wait for Clk_period;
		Addr <=  "0011100001001";
		Trees_din <= x"72ffc808";
		wait for Clk_period;
		Addr <=  "0011100001010";
		Trees_din <= x"51005404";
		wait for Clk_period;
		Addr <=  "0011100001011";
		Trees_din <= x"ffd41c89";
		wait for Clk_period;
		Addr <=  "0011100001100";
		Trees_din <= x"00551c89";
		wait for Clk_period;
		Addr <=  "0011100001101";
		Trees_din <= x"83fe9204";
		wait for Clk_period;
		Addr <=  "0011100001110";
		Trees_din <= x"00071c89";
		wait for Clk_period;
		Addr <=  "0011100001111";
		Trees_din <= x"ff8c1c89";
		wait for Clk_period;
		Addr <=  "0011100010000";
		Trees_din <= x"21ffbc04";
		wait for Clk_period;
		Addr <=  "0011100010001";
		Trees_din <= x"ffea1c89";
		wait for Clk_period;
		Addr <=  "0011100010010";
		Trees_din <= x"00711c89";
		wait for Clk_period;
		Addr <=  "0011100010011";
		Trees_din <= x"a6ff9210";
		wait for Clk_period;
		Addr <=  "0011100010100";
		Trees_din <= x"1cfee308";
		wait for Clk_period;
		Addr <=  "0011100010101";
		Trees_din <= x"ceff4a04";
		wait for Clk_period;
		Addr <=  "0011100010110";
		Trees_din <= x"00591c89";
		wait for Clk_period;
		Addr <=  "0011100010111";
		Trees_din <= x"ffc31c89";
		wait for Clk_period;
		Addr <=  "0011100011000";
		Trees_din <= x"a6fed704";
		wait for Clk_period;
		Addr <=  "0011100011001";
		Trees_din <= x"ffef1c89";
		wait for Clk_period;
		Addr <=  "0011100011010";
		Trees_din <= x"ff751c89";
		wait for Clk_period;
		Addr <=  "0011100011011";
		Trees_din <= x"be001f08";
		wait for Clk_period;
		Addr <=  "0011100011100";
		Trees_din <= x"5a005404";
		wait for Clk_period;
		Addr <=  "0011100011101";
		Trees_din <= x"fff91c89";
		wait for Clk_period;
		Addr <=  "0011100011110";
		Trees_din <= x"ff9f1c89";
		wait for Clk_period;
		Addr <=  "0011100011111";
		Trees_din <= x"ceffc704";
		wait for Clk_period;
		Addr <=  "0011100100000";
		Trees_din <= x"ffff1c89";
		wait for Clk_period;
		Addr <=  "0011100100001";
		Trees_din <= x"008f1c89";
		wait for Clk_period;
		Addr <=  "0011100100010";
		Trees_din <= x"49001064";
		wait for Clk_period;
		Addr <=  "0011100100011";
		Trees_din <= x"28ff2b34";
		wait for Clk_period;
		Addr <=  "0011100100100";
		Trees_din <= x"8a004320";
		wait for Clk_period;
		Addr <=  "0011100100101";
		Trees_din <= x"5a000010";
		wait for Clk_period;
		Addr <=  "0011100100110";
		Trees_din <= x"1cfeff08";
		wait for Clk_period;
		Addr <=  "0011100100111";
		Trees_din <= x"c6ff2504";
		wait for Clk_period;
		Addr <=  "0011100101000";
		Trees_din <= x"000b1da5";
		wait for Clk_period;
		Addr <=  "0011100101001";
		Trees_din <= x"00821da5";
		wait for Clk_period;
		Addr <=  "0011100101010";
		Trees_din <= x"3cff4404";
		wait for Clk_period;
		Addr <=  "0011100101011";
		Trees_din <= x"ff921da5";
		wait for Clk_period;
		Addr <=  "0011100101100";
		Trees_din <= x"001c1da5";
		wait for Clk_period;
		Addr <=  "0011100101101";
		Trees_din <= x"b3fec308";
		wait for Clk_period;
		Addr <=  "0011100101110";
		Trees_din <= x"76ff6604";
		wait for Clk_period;
		Addr <=  "0011100101111";
		Trees_din <= x"005b1da5";
		wait for Clk_period;
		Addr <=  "0011100110000";
		Trees_din <= x"ffb51da5";
		wait for Clk_period;
		Addr <=  "0011100110001";
		Trees_din <= x"2dfe1504";
		wait for Clk_period;
		Addr <=  "0011100110010";
		Trees_din <= x"000b1da5";
		wait for Clk_period;
		Addr <=  "0011100110011";
		Trees_din <= x"ff7d1da5";
		wait for Clk_period;
		Addr <=  "0011100110100";
		Trees_din <= x"faff800c";
		wait for Clk_period;
		Addr <=  "0011100110101";
		Trees_din <= x"1b003f04";
		wait for Clk_period;
		Addr <=  "0011100110110";
		Trees_din <= x"ffab1da5";
		wait for Clk_period;
		Addr <=  "0011100110111";
		Trees_din <= x"f4feba04";
		wait for Clk_period;
		Addr <=  "0011100111000";
		Trees_din <= x"00521da5";
		wait for Clk_period;
		Addr <=  "0011100111001";
		Trees_din <= x"ffe91da5";
		wait for Clk_period;
		Addr <=  "0011100111010";
		Trees_din <= x"81ff8d04";
		wait for Clk_period;
		Addr <=  "0011100111011";
		Trees_din <= x"007d1da5";
		wait for Clk_period;
		Addr <=  "0011100111100";
		Trees_din <= x"fffa1da5";
		wait for Clk_period;
		Addr <=  "0011100111101";
		Trees_din <= x"2fff791c";
		wait for Clk_period;
		Addr <=  "0011100111110";
		Trees_din <= x"e1ffe90c";
		wait for Clk_period;
		Addr <=  "0011100111111";
		Trees_din <= x"ea000008";
		wait for Clk_period;
		Addr <=  "0011101000000";
		Trees_din <= x"43002a04";
		wait for Clk_period;
		Addr <=  "0011101000001";
		Trees_din <= x"ff7a1da5";
		wait for Clk_period;
		Addr <=  "0011101000010";
		Trees_din <= x"00151da5";
		wait for Clk_period;
		Addr <=  "0011101000011";
		Trees_din <= x"004b1da5";
		wait for Clk_period;
		Addr <=  "0011101000100";
		Trees_din <= x"47fffa08";
		wait for Clk_period;
		Addr <=  "0011101000101";
		Trees_din <= x"90fffb04";
		wait for Clk_period;
		Addr <=  "0011101000110";
		Trees_din <= x"ffa01da5";
		wait for Clk_period;
		Addr <=  "0011101000111";
		Trees_din <= x"001b1da5";
		wait for Clk_period;
		Addr <=  "0011101001000";
		Trees_din <= x"16feb604";
		wait for Clk_period;
		Addr <=  "0011101001001";
		Trees_din <= x"ffc31da5";
		wait for Clk_period;
		Addr <=  "0011101001010";
		Trees_din <= x"006c1da5";
		wait for Clk_period;
		Addr <=  "0011101001011";
		Trees_din <= x"4bff3b0c";
		wait for Clk_period;
		Addr <=  "0011101001100";
		Trees_din <= x"abffe404";
		wait for Clk_period;
		Addr <=  "0011101001101";
		Trees_din <= x"ffac1da5";
		wait for Clk_period;
		Addr <=  "0011101001110";
		Trees_din <= x"95ffc804";
		wait for Clk_period;
		Addr <=  "0011101001111";
		Trees_din <= x"006d1da5";
		wait for Clk_period;
		Addr <=  "0011101010000";
		Trees_din <= x"ffbd1da5";
		wait for Clk_period;
		Addr <=  "0011101010001";
		Trees_din <= x"c3ff9804";
		wait for Clk_period;
		Addr <=  "0011101010010";
		Trees_din <= x"003e1da5";
		wait for Clk_period;
		Addr <=  "0011101010011";
		Trees_din <= x"ffa11da5";
		wait for Clk_period;
		Addr <=  "0011101010100";
		Trees_din <= x"e2ff2d20";
		wait for Clk_period;
		Addr <=  "0011101010101";
		Trees_din <= x"11ff880c";
		wait for Clk_period;
		Addr <=  "0011101010110";
		Trees_din <= x"89010608";
		wait for Clk_period;
		Addr <=  "0011101010111";
		Trees_din <= x"84004804";
		wait for Clk_period;
		Addr <=  "0011101011000";
		Trees_din <= x"ff781da5";
		wait for Clk_period;
		Addr <=  "0011101011001";
		Trees_din <= x"001f1da5";
		wait for Clk_period;
		Addr <=  "0011101011010";
		Trees_din <= x"00461da5";
		wait for Clk_period;
		Addr <=  "0011101011011";
		Trees_din <= x"65ff3d0c";
		wait for Clk_period;
		Addr <=  "0011101011100";
		Trees_din <= x"c5ff4708";
		wait for Clk_period;
		Addr <=  "0011101011101";
		Trees_din <= x"f3fea204";
		wait for Clk_period;
		Addr <=  "0011101011110";
		Trees_din <= x"000a1da5";
		wait for Clk_period;
		Addr <=  "0011101011111";
		Trees_din <= x"00871da5";
		wait for Clk_period;
		Addr <=  "0011101100000";
		Trees_din <= x"ffd71da5";
		wait for Clk_period;
		Addr <=  "0011101100001";
		Trees_din <= x"e4fe2904";
		wait for Clk_period;
		Addr <=  "0011101100010";
		Trees_din <= x"00211da5";
		wait for Clk_period;
		Addr <=  "0011101100011";
		Trees_din <= x"ff931da5";
		wait for Clk_period;
		Addr <=  "0011101100100";
		Trees_din <= x"5ffe8c04";
		wait for Clk_period;
		Addr <=  "0011101100101";
		Trees_din <= x"00091da5";
		wait for Clk_period;
		Addr <=  "0011101100110";
		Trees_din <= x"37fee904";
		wait for Clk_period;
		Addr <=  "0011101100111";
		Trees_din <= x"ffe31da5";
		wait for Clk_period;
		Addr <=  "0011101101000";
		Trees_din <= x"ff761da5";
		wait for Clk_period;
		Addr <=  "0011101101001";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0011101101010";
		Trees_din <= x"0fff3138";
		wait for Clk_period;
		Addr <=  "0011101101011";
		Trees_din <= x"f7ff2e14";
		wait for Clk_period;
		Addr <=  "0011101101100";
		Trees_din <= x"dc00b70c";
		wait for Clk_period;
		Addr <=  "0011101101101";
		Trees_din <= x"27007408";
		wait for Clk_period;
		Addr <=  "0011101101110";
		Trees_din <= x"a6feec04";
		wait for Clk_period;
		Addr <=  "0011101101111";
		Trees_din <= x"ffe61e95";
		wait for Clk_period;
		Addr <=  "0011101110000";
		Trees_din <= x"ff7d1e95";
		wait for Clk_period;
		Addr <=  "0011101110001";
		Trees_din <= x"00261e95";
		wait for Clk_period;
		Addr <=  "0011101110010";
		Trees_din <= x"f3feb804";
		wait for Clk_period;
		Addr <=  "0011101110011";
		Trees_din <= x"00081e95";
		wait for Clk_period;
		Addr <=  "0011101110100";
		Trees_din <= x"00641e95";
		wait for Clk_period;
		Addr <=  "0011101110101";
		Trees_din <= x"25ffcb0c";
		wait for Clk_period;
		Addr <=  "0011101110110";
		Trees_din <= x"93feeb04";
		wait for Clk_period;
		Addr <=  "0011101110111";
		Trees_din <= x"002e1e95";
		wait for Clk_period;
		Addr <=  "0011101111000";
		Trees_din <= x"e9febf04";
		wait for Clk_period;
		Addr <=  "0011101111001";
		Trees_din <= x"ffea1e95";
		wait for Clk_period;
		Addr <=  "0011101111010";
		Trees_din <= x"ff9b1e95";
		wait for Clk_period;
		Addr <=  "0011101111011";
		Trees_din <= x"a2ff7208";
		wait for Clk_period;
		Addr <=  "0011101111100";
		Trees_din <= x"7affe504";
		wait for Clk_period;
		Addr <=  "0011101111101";
		Trees_din <= x"ffb71e95";
		wait for Clk_period;
		Addr <=  "0011101111110";
		Trees_din <= x"00341e95";
		wait for Clk_period;
		Addr <=  "0011101111111";
		Trees_din <= x"71ff7a08";
		wait for Clk_period;
		Addr <=  "0011110000000";
		Trees_din <= x"e3fe7a04";
		wait for Clk_period;
		Addr <=  "0011110000001";
		Trees_din <= x"00091e95";
		wait for Clk_period;
		Addr <=  "0011110000010";
		Trees_din <= x"00871e95";
		wait for Clk_period;
		Addr <=  "0011110000011";
		Trees_din <= x"b8ff9c04";
		wait for Clk_period;
		Addr <=  "0011110000100";
		Trees_din <= x"ffa51e95";
		wait for Clk_period;
		Addr <=  "0011110000101";
		Trees_din <= x"00471e95";
		wait for Clk_period;
		Addr <=  "0011110000110";
		Trees_din <= x"30ffb510";
		wait for Clk_period;
		Addr <=  "0011110000111";
		Trees_din <= x"2c00680c";
		wait for Clk_period;
		Addr <=  "0011110001000";
		Trees_din <= x"5cff6904";
		wait for Clk_period;
		Addr <=  "0011110001001";
		Trees_din <= x"fffc1e95";
		wait for Clk_period;
		Addr <=  "0011110001010";
		Trees_din <= x"a5ff9604";
		wait for Clk_period;
		Addr <=  "0011110001011";
		Trees_din <= x"ff721e95";
		wait for Clk_period;
		Addr <=  "0011110001100";
		Trees_din <= x"ffd21e95";
		wait for Clk_period;
		Addr <=  "0011110001101";
		Trees_din <= x"002f1e95";
		wait for Clk_period;
		Addr <=  "0011110001110";
		Trees_din <= x"a9ffb520";
		wait for Clk_period;
		Addr <=  "0011110001111";
		Trees_din <= x"2affdf10";
		wait for Clk_period;
		Addr <=  "0011110010000";
		Trees_din <= x"d3ff4508";
		wait for Clk_period;
		Addr <=  "0011110010001";
		Trees_din <= x"2ffffc04";
		wait for Clk_period;
		Addr <=  "0011110010010";
		Trees_din <= x"ff8d1e95";
		wait for Clk_period;
		Addr <=  "0011110010011";
		Trees_din <= x"00251e95";
		wait for Clk_period;
		Addr <=  "0011110010100";
		Trees_din <= x"aeff4804";
		wait for Clk_period;
		Addr <=  "0011110010101";
		Trees_din <= x"ffc21e95";
		wait for Clk_period;
		Addr <=  "0011110010110";
		Trees_din <= x"00661e95";
		wait for Clk_period;
		Addr <=  "0011110010111";
		Trees_din <= x"49000908";
		wait for Clk_period;
		Addr <=  "0011110011000";
		Trees_din <= x"f7fffb04";
		wait for Clk_period;
		Addr <=  "0011110011001";
		Trees_din <= x"006b1e95";
		wait for Clk_period;
		Addr <=  "0011110011010";
		Trees_din <= x"fff51e95";
		wait for Clk_period;
		Addr <=  "0011110011011";
		Trees_din <= x"3bfebb04";
		wait for Clk_period;
		Addr <=  "0011110011100";
		Trees_din <= x"005f1e95";
		wait for Clk_period;
		Addr <=  "0011110011101";
		Trees_din <= x"ffb61e95";
		wait for Clk_period;
		Addr <=  "0011110011110";
		Trees_din <= x"2e00810c";
		wait for Clk_period;
		Addr <=  "0011110011111";
		Trees_din <= x"9efedc04";
		wait for Clk_period;
		Addr <=  "0011110100000";
		Trees_din <= x"00191e95";
		wait for Clk_period;
		Addr <=  "0011110100001";
		Trees_din <= x"3bfeb404";
		wait for Clk_period;
		Addr <=  "0011110100010";
		Trees_din <= x"ffe91e95";
		wait for Clk_period;
		Addr <=  "0011110100011";
		Trees_din <= x"ff751e95";
		wait for Clk_period;
		Addr <=  "0011110100100";
		Trees_din <= x"00661e95";
		wait for Clk_period;
		Addr <=  "0011110100101";
		Trees_din <= x"8dfe9038";
		wait for Clk_period;
		Addr <=  "0011110100110";
		Trees_din <= x"73ffd510";
		wait for Clk_period;
		Addr <=  "0011110100111";
		Trees_din <= x"3afeb60c";
		wait for Clk_period;
		Addr <=  "0011110101000";
		Trees_din <= x"28ff2a04";
		wait for Clk_period;
		Addr <=  "0011110101001";
		Trees_din <= x"ffa51f81";
		wait for Clk_period;
		Addr <=  "0011110101010";
		Trees_din <= x"04007004";
		wait for Clk_period;
		Addr <=  "0011110101011";
		Trees_din <= x"ffe51f81";
		wait for Clk_period;
		Addr <=  "0011110101100";
		Trees_din <= x"00501f81";
		wait for Clk_period;
		Addr <=  "0011110101101";
		Trees_din <= x"ff7b1f81";
		wait for Clk_period;
		Addr <=  "0011110101110";
		Trees_din <= x"68fe9618";
		wait for Clk_period;
		Addr <=  "0011110101111";
		Trees_din <= x"f7ff4608";
		wait for Clk_period;
		Addr <=  "0011110110000";
		Trees_din <= x"77ff0604";
		wait for Clk_period;
		Addr <=  "0011110110001";
		Trees_din <= x"ffad1f81";
		wait for Clk_period;
		Addr <=  "0011110110010";
		Trees_din <= x"00111f81";
		wait for Clk_period;
		Addr <=  "0011110110011";
		Trees_din <= x"27ffed08";
		wait for Clk_period;
		Addr <=  "0011110110100";
		Trees_din <= x"9bff1004";
		wait for Clk_period;
		Addr <=  "0011110110101";
		Trees_din <= x"002f1f81";
		wait for Clk_period;
		Addr <=  "0011110110110";
		Trees_din <= x"ffc41f81";
		wait for Clk_period;
		Addr <=  "0011110110111";
		Trees_din <= x"7dffe904";
		wait for Clk_period;
		Addr <=  "0011110111000";
		Trees_din <= x"00811f81";
		wait for Clk_period;
		Addr <=  "0011110111001";
		Trees_din <= x"00131f81";
		wait for Clk_period;
		Addr <=  "0011110111010";
		Trees_din <= x"d4ff1804";
		wait for Clk_period;
		Addr <=  "0011110111011";
		Trees_din <= x"ff841f81";
		wait for Clk_period;
		Addr <=  "0011110111100";
		Trees_din <= x"c7fedc08";
		wait for Clk_period;
		Addr <=  "0011110111101";
		Trees_din <= x"7d003804";
		wait for Clk_period;
		Addr <=  "0011110111110";
		Trees_din <= x"ffdd1f81";
		wait for Clk_period;
		Addr <=  "0011110111111";
		Trees_din <= x"00491f81";
		wait for Clk_period;
		Addr <=  "0011111000000";
		Trees_din <= x"ffa21f81";
		wait for Clk_period;
		Addr <=  "0011111000001";
		Trees_din <= x"01fed31c";
		wait for Clk_period;
		Addr <=  "0011111000010";
		Trees_din <= x"e2ff8514";
		wait for Clk_period;
		Addr <=  "0011111000011";
		Trees_din <= x"1aff5110";
		wait for Clk_period;
		Addr <=  "0011111000100";
		Trees_din <= x"8effbd08";
		wait for Clk_period;
		Addr <=  "0011111000101";
		Trees_din <= x"6aff8004";
		wait for Clk_period;
		Addr <=  "0011111000110";
		Trees_din <= x"003a1f81";
		wait for Clk_period;
		Addr <=  "0011111000111";
		Trees_din <= x"ffa21f81";
		wait for Clk_period;
		Addr <=  "0011111001000";
		Trees_din <= x"17ffd404";
		wait for Clk_period;
		Addr <=  "0011111001001";
		Trees_din <= x"000e1f81";
		wait for Clk_period;
		Addr <=  "0011111001010";
		Trees_din <= x"00621f81";
		wait for Clk_period;
		Addr <=  "0011111001011";
		Trees_din <= x"ffbd1f81";
		wait for Clk_period;
		Addr <=  "0011111001100";
		Trees_din <= x"f9ffad04";
		wait for Clk_period;
		Addr <=  "0011111001101";
		Trees_din <= x"ff891f81";
		wait for Clk_period;
		Addr <=  "0011111001110";
		Trees_din <= x"002c1f81";
		wait for Clk_period;
		Addr <=  "0011111001111";
		Trees_din <= x"fcff0e10";
		wait for Clk_period;
		Addr <=  "0011111010000";
		Trees_din <= x"2affac04";
		wait for Clk_period;
		Addr <=  "0011111010001";
		Trees_din <= x"ff991f81";
		wait for Clk_period;
		Addr <=  "0011111010010";
		Trees_din <= x"14fedd04";
		wait for Clk_period;
		Addr <=  "0011111010011";
		Trees_din <= x"ffd21f81";
		wait for Clk_period;
		Addr <=  "0011111010100";
		Trees_din <= x"daffd504";
		wait for Clk_period;
		Addr <=  "0011111010101";
		Trees_din <= x"fff11f81";
		wait for Clk_period;
		Addr <=  "0011111010110";
		Trees_din <= x"00861f81";
		wait for Clk_period;
		Addr <=  "0011111010111";
		Trees_din <= x"a2ff9a08";
		wait for Clk_period;
		Addr <=  "0011111011000";
		Trees_din <= x"08008d04";
		wait for Clk_period;
		Addr <=  "0011111011001";
		Trees_din <= x"ffd11f81";
		wait for Clk_period;
		Addr <=  "0011111011010";
		Trees_din <= x"004f1f81";
		wait for Clk_period;
		Addr <=  "0011111011011";
		Trees_din <= x"4cffe508";
		wait for Clk_period;
		Addr <=  "0011111011100";
		Trees_din <= x"0a00d504";
		wait for Clk_period;
		Addr <=  "0011111011101";
		Trees_din <= x"ff771f81";
		wait for Clk_period;
		Addr <=  "0011111011110";
		Trees_din <= x"ffe21f81";
		wait for Clk_period;
		Addr <=  "0011111011111";
		Trees_din <= x"000f1f81";
		wait for Clk_period;
		Addr <=  "0011111100000";
		Trees_din <= x"a9ff664c";
		wait for Clk_period;
		Addr <=  "0011111100001";
		Trees_din <= x"e2ff2a30";
		wait for Clk_period;
		Addr <=  "0011111100010";
		Trees_din <= x"a0fe8110";
		wait for Clk_period;
		Addr <=  "0011111100011";
		Trees_din <= x"ebff2708";
		wait for Clk_period;
		Addr <=  "0011111100100";
		Trees_din <= x"10ffe304";
		wait for Clk_period;
		Addr <=  "0011111100101";
		Trees_din <= x"ff92208d";
		wait for Clk_period;
		Addr <=  "0011111100110";
		Trees_din <= x"0005208d";
		wait for Clk_period;
		Addr <=  "0011111100111";
		Trees_din <= x"cc001604";
		wait for Clk_period;
		Addr <=  "0011111101000";
		Trees_din <= x"000b208d";
		wait for Clk_period;
		Addr <=  "0011111101001";
		Trees_din <= x"0054208d";
		wait for Clk_period;
		Addr <=  "0011111101010";
		Trees_din <= x"c5ff3d10";
		wait for Clk_period;
		Addr <=  "0011111101011";
		Trees_din <= x"f7fffb08";
		wait for Clk_period;
		Addr <=  "0011111101100";
		Trees_din <= x"f1ff5804";
		wait for Clk_period;
		Addr <=  "0011111101101";
		Trees_din <= x"0012208d";
		wait for Clk_period;
		Addr <=  "0011111101110";
		Trees_din <= x"0081208d";
		wait for Clk_period;
		Addr <=  "0011111101111";
		Trees_din <= x"0fff2f04";
		wait for Clk_period;
		Addr <=  "0011111110000";
		Trees_din <= x"0051208d";
		wait for Clk_period;
		Addr <=  "0011111110001";
		Trees_din <= x"ffc5208d";
		wait for Clk_period;
		Addr <=  "0011111110010";
		Trees_din <= x"d6005208";
		wait for Clk_period;
		Addr <=  "0011111110011";
		Trees_din <= x"c6feb004";
		wait for Clk_period;
		Addr <=  "0011111110100";
		Trees_din <= x"0022208d";
		wait for Clk_period;
		Addr <=  "0011111110101";
		Trees_din <= x"ff95208d";
		wait for Clk_period;
		Addr <=  "0011111110110";
		Trees_din <= x"5c004104";
		wait for Clk_period;
		Addr <=  "0011111110111";
		Trees_din <= x"005d208d";
		wait for Clk_period;
		Addr <=  "0011111111000";
		Trees_din <= x"ffe8208d";
		wait for Clk_period;
		Addr <=  "0011111111001";
		Trees_din <= x"5a003910";
		wait for Clk_period;
		Addr <=  "0011111111010";
		Trees_din <= x"0fffa10c";
		wait for Clk_period;
		Addr <=  "0011111111011";
		Trees_din <= x"8dfec904";
		wait for Clk_period;
		Addr <=  "0011111111100";
		Trees_din <= x"ffec208d";
		wait for Clk_period;
		Addr <=  "0011111111101";
		Trees_din <= x"d4ff5304";
		wait for Clk_period;
		Addr <=  "0011111111110";
		Trees_din <= x"0077208d";
		wait for Clk_period;
		Addr <=  "0011111111111";
		Trees_din <= x"0013208d";
		wait for Clk_period;
		Addr <=  "0100000000000";
		Trees_din <= x"ffae208d";
		wait for Clk_period;
		Addr <=  "0100000000001";
		Trees_din <= x"58ffa108";
		wait for Clk_period;
		Addr <=  "0100000000010";
		Trees_din <= x"55008004";
		wait for Clk_period;
		Addr <=  "0100000000011";
		Trees_din <= x"ff7c208d";
		wait for Clk_period;
		Addr <=  "0100000000100";
		Trees_din <= x"fffd208d";
		wait for Clk_period;
		Addr <=  "0100000000101";
		Trees_din <= x"001c208d";
		wait for Clk_period;
		Addr <=  "0100000000110";
		Trees_din <= x"0a002d10";
		wait for Clk_period;
		Addr <=  "0100000000111";
		Trees_din <= x"13019d08";
		wait for Clk_period;
		Addr <=  "0100000001000";
		Trees_din <= x"74ff6f04";
		wait for Clk_period;
		Addr <=  "0100000001001";
		Trees_din <= x"002f208d";
		wait for Clk_period;
		Addr <=  "0100000001010";
		Trees_din <= x"ff76208d";
		wait for Clk_period;
		Addr <=  "0100000001011";
		Trees_din <= x"11ffaf04";
		wait for Clk_period;
		Addr <=  "0100000001100";
		Trees_din <= x"ffe1208d";
		wait for Clk_period;
		Addr <=  "0100000001101";
		Trees_din <= x"0055208d";
		wait for Clk_period;
		Addr <=  "0100000001110";
		Trees_din <= x"e7ff9d1c";
		wait for Clk_period;
		Addr <=  "0100000001111";
		Trees_din <= x"1eff9010";
		wait for Clk_period;
		Addr <=  "0100000010000";
		Trees_din <= x"59ff8b08";
		wait for Clk_period;
		Addr <=  "0100000010001";
		Trees_din <= x"e4fe1904";
		wait for Clk_period;
		Addr <=  "0100000010010";
		Trees_din <= x"fffd208d";
		wait for Clk_period;
		Addr <=  "0100000010011";
		Trees_din <= x"ff89208d";
		wait for Clk_period;
		Addr <=  "0100000010100";
		Trees_din <= x"fcff1304";
		wait for Clk_period;
		Addr <=  "0100000010101";
		Trees_din <= x"0060208d";
		wait for Clk_period;
		Addr <=  "0100000010110";
		Trees_din <= x"ffd8208d";
		wait for Clk_period;
		Addr <=  "0100000010111";
		Trees_din <= x"07002404";
		wait for Clk_period;
		Addr <=  "0100000011000";
		Trees_din <= x"ffbe208d";
		wait for Clk_period;
		Addr <=  "0100000011001";
		Trees_din <= x"17ffc404";
		wait for Clk_period;
		Addr <=  "0100000011010";
		Trees_din <= x"ffe4208d";
		wait for Clk_period;
		Addr <=  "0100000011011";
		Trees_din <= x"005f208d";
		wait for Clk_period;
		Addr <=  "0100000011100";
		Trees_din <= x"e100cb0c";
		wait for Clk_period;
		Addr <=  "0100000011101";
		Trees_din <= x"fb002408";
		wait for Clk_period;
		Addr <=  "0100000011110";
		Trees_din <= x"81ff3004";
		wait for Clk_period;
		Addr <=  "0100000011111";
		Trees_din <= x"ffe3208d";
		wait for Clk_period;
		Addr <=  "0100000100000";
		Trees_din <= x"ff7b208d";
		wait for Clk_period;
		Addr <=  "0100000100001";
		Trees_din <= x"0026208d";
		wait for Clk_period;
		Addr <=  "0100000100010";
		Trees_din <= x"003a208d";
		wait for Clk_period;
		Addr <=  "0100000100011";
		Trees_din <= x"2cff6a24";
		wait for Clk_period;
		Addr <=  "0100000100100";
		Trees_din <= x"b7ff0c08";
		wait for Clk_period;
		Addr <=  "0100000100101";
		Trees_din <= x"fdff2304";
		wait for Clk_period;
		Addr <=  "0100000100110";
		Trees_din <= x"00592169";
		wait for Clk_period;
		Addr <=  "0100000100111";
		Trees_din <= x"ffd92169";
		wait for Clk_period;
		Addr <=  "0100000101000";
		Trees_din <= x"c5ff3014";
		wait for Clk_period;
		Addr <=  "0100000101001";
		Trees_din <= x"0eff200c";
		wait for Clk_period;
		Addr <=  "0100000101010";
		Trees_din <= x"01fe2804";
		wait for Clk_period;
		Addr <=  "0100000101011";
		Trees_din <= x"002b2169";
		wait for Clk_period;
		Addr <=  "0100000101100";
		Trees_din <= x"eaffce04";
		wait for Clk_period;
		Addr <=  "0100000101101";
		Trees_din <= x"ff872169";
		wait for Clk_period;
		Addr <=  "0100000101110";
		Trees_din <= x"00052169";
		wait for Clk_period;
		Addr <=  "0100000101111";
		Trees_din <= x"00ff9b04";
		wait for Clk_period;
		Addr <=  "0100000110000";
		Trees_din <= x"ffdb2169";
		wait for Clk_period;
		Addr <=  "0100000110001";
		Trees_din <= x"00582169";
		wait for Clk_period;
		Addr <=  "0100000110010";
		Trees_din <= x"e1007d04";
		wait for Clk_period;
		Addr <=  "0100000110011";
		Trees_din <= x"ff7a2169";
		wait for Clk_period;
		Addr <=  "0100000110100";
		Trees_din <= x"fffd2169";
		wait for Clk_period;
		Addr <=  "0100000110101";
		Trees_din <= x"73ffc620";
		wait for Clk_period;
		Addr <=  "0100000110110";
		Trees_din <= x"0dff6214";
		wait for Clk_period;
		Addr <=  "0100000110111";
		Trees_din <= x"c7feff0c";
		wait for Clk_period;
		Addr <=  "0100000111000";
		Trees_din <= x"4eff0c04";
		wait for Clk_period;
		Addr <=  "0100000111001";
		Trees_din <= x"ffc32169";
		wait for Clk_period;
		Addr <=  "0100000111010";
		Trees_din <= x"c1fe8904";
		wait for Clk_period;
		Addr <=  "0100000111011";
		Trees_din <= x"ffe12169";
		wait for Clk_period;
		Addr <=  "0100000111100";
		Trees_din <= x"00582169";
		wait for Clk_period;
		Addr <=  "0100000111101";
		Trees_din <= x"0ffefa04";
		wait for Clk_period;
		Addr <=  "0100000111110";
		Trees_din <= x"00132169";
		wait for Clk_period;
		Addr <=  "0100000111111";
		Trees_din <= x"ff972169";
		wait for Clk_period;
		Addr <=  "0100001000000";
		Trees_din <= x"b4ffa808";
		wait for Clk_period;
		Addr <=  "0100001000001";
		Trees_din <= x"d8fff804";
		wait for Clk_period;
		Addr <=  "0100001000010";
		Trees_din <= x"ffdc2169";
		wait for Clk_period;
		Addr <=  "0100001000011";
		Trees_din <= x"ff7e2169";
		wait for Clk_period;
		Addr <=  "0100001000100";
		Trees_din <= x"000d2169";
		wait for Clk_period;
		Addr <=  "0100001000101";
		Trees_din <= x"14ff6d20";
		wait for Clk_period;
		Addr <=  "0100001000110";
		Trees_din <= x"5cffbf10";
		wait for Clk_period;
		Addr <=  "0100001000111";
		Trees_din <= x"2affbc08";
		wait for Clk_period;
		Addr <=  "0100001001000";
		Trees_din <= x"50ff1f04";
		wait for Clk_period;
		Addr <=  "0100001001001";
		Trees_din <= x"00332169";
		wait for Clk_period;
		Addr <=  "0100001001010";
		Trees_din <= x"ffaa2169";
		wait for Clk_period;
		Addr <=  "0100001001011";
		Trees_din <= x"96ff2a04";
		wait for Clk_period;
		Addr <=  "0100001001100";
		Trees_din <= x"00052169";
		wait for Clk_period;
		Addr <=  "0100001001101";
		Trees_din <= x"007b2169";
		wait for Clk_period;
		Addr <=  "0100001001110";
		Trees_din <= x"19ff4908";
		wait for Clk_period;
		Addr <=  "0100001001111";
		Trees_din <= x"36ffc604";
		wait for Clk_period;
		Addr <=  "0100001010000";
		Trees_din <= x"00412169";
		wait for Clk_period;
		Addr <=  "0100001010001";
		Trees_din <= x"ffb42169";
		wait for Clk_period;
		Addr <=  "0100001010010";
		Trees_din <= x"0a00c604";
		wait for Clk_period;
		Addr <=  "0100001010011";
		Trees_din <= x"ffa92169";
		wait for Clk_period;
		Addr <=  "0100001010100";
		Trees_din <= x"00282169";
		wait for Clk_period;
		Addr <=  "0100001010101";
		Trees_din <= x"7fffb204";
		wait for Clk_period;
		Addr <=  "0100001010110";
		Trees_din <= x"ff902169";
		wait for Clk_period;
		Addr <=  "0100001010111";
		Trees_din <= x"39ff7404";
		wait for Clk_period;
		Addr <=  "0100001011000";
		Trees_din <= x"00602169";
		wait for Clk_period;
		Addr <=  "0100001011001";
		Trees_din <= x"ffd42169";
		wait for Clk_period;
		Addr <=  "0100001011010";
		Trees_din <= x"aaff7344";
		wait for Clk_period;
		Addr <=  "0100001011011";
		Trees_din <= x"b4fe9a20";
		wait for Clk_period;
		Addr <=  "0100001011100";
		Trees_din <= x"bbff5a10";
		wait for Clk_period;
		Addr <=  "0100001011101";
		Trees_din <= x"a1fec304";
		wait for Clk_period;
		Addr <=  "0100001011110";
		Trees_din <= x"ff9c2265";
		wait for Clk_period;
		Addr <=  "0100001011111";
		Trees_din <= x"c8001f04";
		wait for Clk_period;
		Addr <=  "0100001100000";
		Trees_din <= x"ffd12265";
		wait for Clk_period;
		Addr <=  "0100001100001";
		Trees_din <= x"9fff6104";
		wait for Clk_period;
		Addr <=  "0100001100010";
		Trees_din <= x"00012265";
		wait for Clk_period;
		Addr <=  "0100001100011";
		Trees_din <= x"00562265";
		wait for Clk_period;
		Addr <=  "0100001100100";
		Trees_din <= x"33feb504";
		wait for Clk_period;
		Addr <=  "0100001100101";
		Trees_din <= x"ffc92265";
		wait for Clk_period;
		Addr <=  "0100001100110";
		Trees_din <= x"ceffd908";
		wait for Clk_period;
		Addr <=  "0100001100111";
		Trees_din <= x"f7ff2e04";
		wait for Clk_period;
		Addr <=  "0100001101000";
		Trees_din <= x"00162265";
		wait for Clk_period;
		Addr <=  "0100001101001";
		Trees_din <= x"007c2265";
		wait for Clk_period;
		Addr <=  "0100001101010";
		Trees_din <= x"ffe92265";
		wait for Clk_period;
		Addr <=  "0100001101011";
		Trees_din <= x"0cfe2e10";
		wait for Clk_period;
		Addr <=  "0100001101100";
		Trees_din <= x"daffbc04";
		wait for Clk_period;
		Addr <=  "0100001101101";
		Trees_din <= x"ffac2265";
		wait for Clk_period;
		Addr <=  "0100001101110";
		Trees_din <= x"1bffb604";
		wait for Clk_period;
		Addr <=  "0100001101111";
		Trees_din <= x"ffd42265";
		wait for Clk_period;
		Addr <=  "0100001110000";
		Trees_din <= x"afffd704";
		wait for Clk_period;
		Addr <=  "0100001110001";
		Trees_din <= x"000a2265";
		wait for Clk_period;
		Addr <=  "0100001110010";
		Trees_din <= x"006d2265";
		wait for Clk_period;
		Addr <=  "0100001110011";
		Trees_din <= x"faffa508";
		wait for Clk_period;
		Addr <=  "0100001110100";
		Trees_din <= x"5e003704";
		wait for Clk_period;
		Addr <=  "0100001110101";
		Trees_din <= x"ff762265";
		wait for Clk_period;
		Addr <=  "0100001110110";
		Trees_din <= x"ffd22265";
		wait for Clk_period;
		Addr <=  "0100001110111";
		Trees_din <= x"c7fe8304";
		wait for Clk_period;
		Addr <=  "0100001111000";
		Trees_din <= x"002a2265";
		wait for Clk_period;
		Addr <=  "0100001111001";
		Trees_din <= x"8e004004";
		wait for Clk_period;
		Addr <=  "0100001111010";
		Trees_din <= x"ff9a2265";
		wait for Clk_period;
		Addr <=  "0100001111011";
		Trees_din <= x"fff72265";
		wait for Clk_period;
		Addr <=  "0100001111100";
		Trees_din <= x"ee006d34";
		wait for Clk_period;
		Addr <=  "0100001111101";
		Trees_din <= x"e2ff231c";
		wait for Clk_period;
		Addr <=  "0100001111110";
		Trees_din <= x"a9ff720c";
		wait for Clk_period;
		Addr <=  "0100001111111";
		Trees_din <= x"f4fe6b04";
		wait for Clk_period;
		Addr <=  "0100010000000";
		Trees_din <= x"ffd02265";
		wait for Clk_period;
		Addr <=  "0100010000001";
		Trees_din <= x"ebfed904";
		wait for Clk_period;
		Addr <=  "0100010000010";
		Trees_din <= x"00082265";
		wait for Clk_period;
		Addr <=  "0100010000011";
		Trees_din <= x"00752265";
		wait for Clk_period;
		Addr <=  "0100010000100";
		Trees_din <= x"8a004308";
		wait for Clk_period;
		Addr <=  "0100010000101";
		Trees_din <= x"fbffff04";
		wait for Clk_period;
		Addr <=  "0100010000110";
		Trees_din <= x"ffa82265";
		wait for Clk_period;
		Addr <=  "0100010000111";
		Trees_din <= x"002b2265";
		wait for Clk_period;
		Addr <=  "0100010001000";
		Trees_din <= x"77ff8c04";
		wait for Clk_period;
		Addr <=  "0100010001001";
		Trees_din <= x"000c2265";
		wait for Clk_period;
		Addr <=  "0100010001010";
		Trees_din <= x"005e2265";
		wait for Clk_period;
		Addr <=  "0100010001011";
		Trees_din <= x"43ff4108";
		wait for Clk_period;
		Addr <=  "0100010001100";
		Trees_din <= x"7fffce04";
		wait for Clk_period;
		Addr <=  "0100010001101";
		Trees_din <= x"ff8d2265";
		wait for Clk_period;
		Addr <=  "0100010001110";
		Trees_din <= x"fff52265";
		wait for Clk_period;
		Addr <=  "0100010001111";
		Trees_din <= x"49001008";
		wait for Clk_period;
		Addr <=  "0100010010000";
		Trees_din <= x"2cff7104";
		wait for Clk_period;
		Addr <=  "0100010010001";
		Trees_din <= x"ffbb2265";
		wait for Clk_period;
		Addr <=  "0100010010010";
		Trees_din <= x"003c2265";
		wait for Clk_period;
		Addr <=  "0100010010011";
		Trees_din <= x"66fff604";
		wait for Clk_period;
		Addr <=  "0100010010100";
		Trees_din <= x"ff9b2265";
		wait for Clk_period;
		Addr <=  "0100010010101";
		Trees_din <= x"fffb2265";
		wait for Clk_period;
		Addr <=  "0100010010110";
		Trees_din <= x"a7001804";
		wait for Clk_period;
		Addr <=  "0100010010111";
		Trees_din <= x"ff942265";
		wait for Clk_period;
		Addr <=  "0100010011000";
		Trees_din <= x"fffc2265";
		wait for Clk_period;
		Addr <=  "0100010011001";
		Trees_din <= x"9cff9444";
		wait for Clk_period;
		Addr <=  "0100010011010";
		Trees_din <= x"c7fee62c";
		wait for Clk_period;
		Addr <=  "0100010011011";
		Trees_din <= x"90ff9714";
		wait for Clk_period;
		Addr <=  "0100010011100";
		Trees_din <= x"43ffde0c";
		wait for Clk_period;
		Addr <=  "0100010011101";
		Trees_din <= x"ccff0604";
		wait for Clk_period;
		Addr <=  "0100010011110";
		Trees_din <= x"002c2361";
		wait for Clk_period;
		Addr <=  "0100010011111";
		Trees_din <= x"49ffa004";
		wait for Clk_period;
		Addr <=  "0100010100000";
		Trees_din <= x"fffb2361";
		wait for Clk_period;
		Addr <=  "0100010100001";
		Trees_din <= x"ff872361";
		wait for Clk_period;
		Addr <=  "0100010100010";
		Trees_din <= x"46feaa04";
		wait for Clk_period;
		Addr <=  "0100010100011";
		Trees_din <= x"005a2361";
		wait for Clk_period;
		Addr <=  "0100010100100";
		Trees_din <= x"00012361";
		wait for Clk_period;
		Addr <=  "0100010100101";
		Trees_din <= x"faff6c0c";
		wait for Clk_period;
		Addr <=  "0100010100110";
		Trees_din <= x"8e003304";
		wait for Clk_period;
		Addr <=  "0100010100111";
		Trees_din <= x"ffa62361";
		wait for Clk_period;
		Addr <=  "0100010101000";
		Trees_din <= x"ccffea04";
		wait for Clk_period;
		Addr <=  "0100010101001";
		Trees_din <= x"fff22361";
		wait for Clk_period;
		Addr <=  "0100010101010";
		Trees_din <= x"00512361";
		wait for Clk_period;
		Addr <=  "0100010101011";
		Trees_din <= x"8aff8a04";
		wait for Clk_period;
		Addr <=  "0100010101100";
		Trees_din <= x"fff32361";
		wait for Clk_period;
		Addr <=  "0100010101101";
		Trees_din <= x"adffbd04";
		wait for Clk_period;
		Addr <=  "0100010101110";
		Trees_din <= x"006f2361";
		wait for Clk_period;
		Addr <=  "0100010101111";
		Trees_din <= x"00002361";
		wait for Clk_period;
		Addr <=  "0100010110000";
		Trees_din <= x"2ffff410";
		wait for Clk_period;
		Addr <=  "0100010110001";
		Trees_din <= x"50fef008";
		wait for Clk_period;
		Addr <=  "0100010110010";
		Trees_din <= x"b2ffec04";
		wait for Clk_period;
		Addr <=  "0100010110011";
		Trees_din <= x"ffda2361";
		wait for Clk_period;
		Addr <=  "0100010110100";
		Trees_din <= x"00392361";
		wait for Clk_period;
		Addr <=  "0100010110101";
		Trees_din <= x"e4fe1904";
		wait for Clk_period;
		Addr <=  "0100010110110";
		Trees_din <= x"ffec2361";
		wait for Clk_period;
		Addr <=  "0100010110111";
		Trees_din <= x"ff792361";
		wait for Clk_period;
		Addr <=  "0100010111000";
		Trees_din <= x"db005a04";
		wait for Clk_period;
		Addr <=  "0100010111001";
		Trees_din <= x"ffcb2361";
		wait for Clk_period;
		Addr <=  "0100010111010";
		Trees_din <= x"00432361";
		wait for Clk_period;
		Addr <=  "0100010111011";
		Trees_din <= x"2cff3b08";
		wait for Clk_period;
		Addr <=  "0100010111100";
		Trees_din <= x"4effb504";
		wait for Clk_period;
		Addr <=  "0100010111101";
		Trees_din <= x"ff9a2361";
		wait for Clk_period;
		Addr <=  "0100010111110";
		Trees_din <= x"fffc2361";
		wait for Clk_period;
		Addr <=  "0100010111111";
		Trees_din <= x"c3ffe318";
		wait for Clk_period;
		Addr <=  "0100011000000";
		Trees_din <= x"2fff5f0c";
		wait for Clk_period;
		Addr <=  "0100011000001";
		Trees_din <= x"d6006404";
		wait for Clk_period;
		Addr <=  "0100011000010";
		Trees_din <= x"ffaa2361";
		wait for Clk_period;
		Addr <=  "0100011000011";
		Trees_din <= x"f1ffcb04";
		wait for Clk_period;
		Addr <=  "0100011000100";
		Trees_din <= x"ffdd2361";
		wait for Clk_period;
		Addr <=  "0100011000101";
		Trees_din <= x"005d2361";
		wait for Clk_period;
		Addr <=  "0100011000110";
		Trees_din <= x"9c002108";
		wait for Clk_period;
		Addr <=  "0100011000111";
		Trees_din <= x"de005c04";
		wait for Clk_period;
		Addr <=  "0100011001000";
		Trees_din <= x"00662361";
		wait for Clk_period;
		Addr <=  "0100011001001";
		Trees_din <= x"fff72361";
		wait for Clk_period;
		Addr <=  "0100011001010";
		Trees_din <= x"ffee2361";
		wait for Clk_period;
		Addr <=  "0100011001011";
		Trees_din <= x"55004b10";
		wait for Clk_period;
		Addr <=  "0100011001100";
		Trees_din <= x"21ff8508";
		wait for Clk_period;
		Addr <=  "0100011001101";
		Trees_din <= x"39ff7a04";
		wait for Clk_period;
		Addr <=  "0100011001110";
		Trees_din <= x"00372361";
		wait for Clk_period;
		Addr <=  "0100011001111";
		Trees_din <= x"ffbf2361";
		wait for Clk_period;
		Addr <=  "0100011010000";
		Trees_din <= x"b4feae04";
		wait for Clk_period;
		Addr <=  "0100011010001";
		Trees_din <= x"ffef2361";
		wait for Clk_period;
		Addr <=  "0100011010010";
		Trees_din <= x"ff8a2361";
		wait for Clk_period;
		Addr <=  "0100011010011";
		Trees_din <= x"5fff3e04";
		wait for Clk_period;
		Addr <=  "0100011010100";
		Trees_din <= x"ffe12361";
		wait for Clk_period;
		Addr <=  "0100011010101";
		Trees_din <= x"c4ff2304";
		wait for Clk_period;
		Addr <=  "0100011010110";
		Trees_din <= x"00112361";
		wait for Clk_period;
		Addr <=  "0100011010111";
		Trees_din <= x"006e2361";
		wait for Clk_period;
		Addr <=  "0100011011000";
		Trees_din <= x"30004d54";
		wait for Clk_period;
		Addr <=  "0100011011001";
		Trees_din <= x"89007f38";
		wait for Clk_period;
		Addr <=  "0100011011010";
		Trees_din <= x"4eff9918";
		wait for Clk_period;
		Addr <=  "0100011011011";
		Trees_din <= x"ccff0308";
		wait for Clk_period;
		Addr <=  "0100011011100";
		Trees_din <= x"f9fecc04";
		wait for Clk_period;
		Addr <=  "0100011011101";
		Trees_din <= x"00522435";
		wait for Clk_period;
		Addr <=  "0100011011110";
		Trees_din <= x"ffdb2435";
		wait for Clk_period;
		Addr <=  "0100011011111";
		Trees_din <= x"51ff4908";
		wait for Clk_period;
		Addr <=  "0100011100000";
		Trees_din <= x"38ffa004";
		wait for Clk_period;
		Addr <=  "0100011100001";
		Trees_din <= x"ffab2435";
		wait for Clk_period;
		Addr <=  "0100011100010";
		Trees_din <= x"00412435";
		wait for Clk_period;
		Addr <=  "0100011100011";
		Trees_din <= x"f800e904";
		wait for Clk_period;
		Addr <=  "0100011100100";
		Trees_din <= x"ff902435";
		wait for Clk_period;
		Addr <=  "0100011100101";
		Trees_din <= x"00192435";
		wait for Clk_period;
		Addr <=  "0100011100110";
		Trees_din <= x"7fff9610";
		wait for Clk_period;
		Addr <=  "0100011100111";
		Trees_din <= x"89002f08";
		wait for Clk_period;
		Addr <=  "0100011101000";
		Trees_din <= x"5c00c004";
		wait for Clk_period;
		Addr <=  "0100011101001";
		Trees_din <= x"ff972435";
		wait for Clk_period;
		Addr <=  "0100011101010";
		Trees_din <= x"00312435";
		wait for Clk_period;
		Addr <=  "0100011101011";
		Trees_din <= x"2200ac04";
		wait for Clk_period;
		Addr <=  "0100011101100";
		Trees_din <= x"ffe82435";
		wait for Clk_period;
		Addr <=  "0100011101101";
		Trees_din <= x"004e2435";
		wait for Clk_period;
		Addr <=  "0100011101110";
		Trees_din <= x"05003e08";
		wait for Clk_period;
		Addr <=  "0100011101111";
		Trees_din <= x"26000f04";
		wait for Clk_period;
		Addr <=  "0100011110000";
		Trees_din <= x"00362435";
		wait for Clk_period;
		Addr <=  "0100011110001";
		Trees_din <= x"ffb42435";
		wait for Clk_period;
		Addr <=  "0100011110010";
		Trees_din <= x"16ff3104";
		wait for Clk_period;
		Addr <=  "0100011110011";
		Trees_din <= x"006c2435";
		wait for Clk_period;
		Addr <=  "0100011110100";
		Trees_din <= x"ffe02435";
		wait for Clk_period;
		Addr <=  "0100011110101";
		Trees_din <= x"8effcd08";
		wait for Clk_period;
		Addr <=  "0100011110110";
		Trees_din <= x"dcfff004";
		wait for Clk_period;
		Addr <=  "0100011110111";
		Trees_din <= x"ffa42435";
		wait for Clk_period;
		Addr <=  "0100011111000";
		Trees_din <= x"00072435";
		wait for Clk_period;
		Addr <=  "0100011111001";
		Trees_din <= x"1f00c00c";
		wait for Clk_period;
		Addr <=  "0100011111010";
		Trees_din <= x"1eff4d04";
		wait for Clk_period;
		Addr <=  "0100011111011";
		Trees_din <= x"fff92435";
		wait for Clk_period;
		Addr <=  "0100011111100";
		Trees_din <= x"5effc604";
		wait for Clk_period;
		Addr <=  "0100011111101";
		Trees_din <= x"00162435";
		wait for Clk_period;
		Addr <=  "0100011111110";
		Trees_din <= x"00702435";
		wait for Clk_period;
		Addr <=  "0100011111111";
		Trees_din <= x"55fffe04";
		wait for Clk_period;
		Addr <=  "0100100000000";
		Trees_din <= x"001b2435";
		wait for Clk_period;
		Addr <=  "0100100000001";
		Trees_din <= x"ffb12435";
		wait for Clk_period;
		Addr <=  "0100100000010";
		Trees_din <= x"17ffd008";
		wait for Clk_period;
		Addr <=  "0100100000011";
		Trees_din <= x"88006904";
		wait for Clk_period;
		Addr <=  "0100100000100";
		Trees_din <= x"ffad2435";
		wait for Clk_period;
		Addr <=  "0100100000101";
		Trees_din <= x"00232435";
		wait for Clk_period;
		Addr <=  "0100100000110";
		Trees_din <= x"1f00610c";
		wait for Clk_period;
		Addr <=  "0100100000111";
		Trees_din <= x"39ffcf08";
		wait for Clk_period;
		Addr <=  "0100100001000";
		Trees_din <= x"90ff9c04";
		wait for Clk_period;
		Addr <=  "0100100001001";
		Trees_din <= x"001d2435";
		wait for Clk_period;
		Addr <=  "0100100001010";
		Trees_din <= x"007b2435";
		wait for Clk_period;
		Addr <=  "0100100001011";
		Trees_din <= x"00022435";
		wait for Clk_period;
		Addr <=  "0100100001100";
		Trees_din <= x"ffef2435";
		wait for Clk_period;
		Addr <=  "0100100001101";
		Trees_din <= x"8dfea138";
		wait for Clk_period;
		Addr <=  "0100100001110";
		Trees_din <= x"e6ff9f24";
		wait for Clk_period;
		Addr <=  "0100100001111";
		Trees_din <= x"d000d514";
		wait for Clk_period;
		Addr <=  "0100100010000";
		Trees_din <= x"85ff4508";
		wait for Clk_period;
		Addr <=  "0100100010001";
		Trees_din <= x"fcff1904";
		wait for Clk_period;
		Addr <=  "0100100010010";
		Trees_din <= x"004c2531";
		wait for Clk_period;
		Addr <=  "0100100010011";
		Trees_din <= x"ffdd2531";
		wait for Clk_period;
		Addr <=  "0100100010100";
		Trees_din <= x"a4ff2704";
		wait for Clk_period;
		Addr <=  "0100100010101";
		Trees_din <= x"000f2531";
		wait for Clk_period;
		Addr <=  "0100100010110";
		Trees_din <= x"d8002204";
		wait for Clk_period;
		Addr <=  "0100100010111";
		Trees_din <= x"fff02531";
		wait for Clk_period;
		Addr <=  "0100100011000";
		Trees_din <= x"ff8c2531";
		wait for Clk_period;
		Addr <=  "0100100011001";
		Trees_din <= x"96ff1c04";
		wait for Clk_period;
		Addr <=  "0100100011010";
		Trees_din <= x"ffe02531";
		wait for Clk_period;
		Addr <=  "0100100011011";
		Trees_din <= x"afff7e04";
		wait for Clk_period;
		Addr <=  "0100100011100";
		Trees_din <= x"00042531";
		wait for Clk_period;
		Addr <=  "0100100011101";
		Trees_din <= x"0dff5404";
		wait for Clk_period;
		Addr <=  "0100100011110";
		Trees_din <= x"006c2531";
		wait for Clk_period;
		Addr <=  "0100100011111";
		Trees_din <= x"00172531";
		wait for Clk_period;
		Addr <=  "0100100100000";
		Trees_din <= x"ccff560c";
		wait for Clk_period;
		Addr <=  "0100100100001";
		Trees_din <= x"faff6604";
		wait for Clk_period;
		Addr <=  "0100100100010";
		Trees_din <= x"ffbd2531";
		wait for Clk_period;
		Addr <=  "0100100100011";
		Trees_din <= x"27002004";
		wait for Clk_period;
		Addr <=  "0100100100100";
		Trees_din <= x"fff72531";
		wait for Clk_period;
		Addr <=  "0100100100101";
		Trees_din <= x"00512531";
		wait for Clk_period;
		Addr <=  "0100100100110";
		Trees_din <= x"0a00c804";
		wait for Clk_period;
		Addr <=  "0100100100111";
		Trees_din <= x"ff7f2531";
		wait for Clk_period;
		Addr <=  "0100100101000";
		Trees_din <= x"ffed2531";
		wait for Clk_period;
		Addr <=  "0100100101001";
		Trees_din <= x"c7fee624";
		wait for Clk_period;
		Addr <=  "0100100101010";
		Trees_din <= x"a9ff6610";
		wait for Clk_period;
		Addr <=  "0100100101011";
		Trees_din <= x"3100640c";
		wait for Clk_period;
		Addr <=  "0100100101100";
		Trees_din <= x"0bff8d04";
		wait for Clk_period;
		Addr <=  "0100100101101";
		Trees_din <= x"00022531";
		wait for Clk_period;
		Addr <=  "0100100101110";
		Trees_din <= x"c1fe7904";
		wait for Clk_period;
		Addr <=  "0100100101111";
		Trees_din <= x"00112531";
		wait for Clk_period;
		Addr <=  "0100100110000";
		Trees_din <= x"00712531";
		wait for Clk_period;
		Addr <=  "0100100110001";
		Trees_din <= x"fff02531";
		wait for Clk_period;
		Addr <=  "0100100110010";
		Trees_din <= x"e7ff9d10";
		wait for Clk_period;
		Addr <=  "0100100110011";
		Trees_din <= x"faff8b08";
		wait for Clk_period;
		Addr <=  "0100100110100";
		Trees_din <= x"23002004";
		wait for Clk_period;
		Addr <=  "0100100110101";
		Trees_din <= x"ffad2531";
		wait for Clk_period;
		Addr <=  "0100100110110";
		Trees_din <= x"002e2531";
		wait for Clk_period;
		Addr <=  "0100100110111";
		Trees_din <= x"11ff7704";
		wait for Clk_period;
		Addr <=  "0100100111000";
		Trees_din <= x"000b2531";
		wait for Clk_period;
		Addr <=  "0100100111001";
		Trees_din <= x"005b2531";
		wait for Clk_period;
		Addr <=  "0100100111010";
		Trees_din <= x"ffad2531";
		wait for Clk_period;
		Addr <=  "0100100111011";
		Trees_din <= x"db001f0c";
		wait for Clk_period;
		Addr <=  "0100100111100";
		Trees_din <= x"ccff0e04";
		wait for Clk_period;
		Addr <=  "0100100111101";
		Trees_din <= x"00242531";
		wait for Clk_period;
		Addr <=  "0100100111110";
		Trees_din <= x"0fff0c04";
		wait for Clk_period;
		Addr <=  "0100100111111";
		Trees_din <= x"fff82531";
		wait for Clk_period;
		Addr <=  "0100101000000";
		Trees_din <= x"ff852531";
		wait for Clk_period;
		Addr <=  "0100101000001";
		Trees_din <= x"66ffac08";
		wait for Clk_period;
		Addr <=  "0100101000010";
		Trees_din <= x"c3ff9304";
		wait for Clk_period;
		Addr <=  "0100101000011";
		Trees_din <= x"00192531";
		wait for Clk_period;
		Addr <=  "0100101000100";
		Trees_din <= x"ffa02531";
		wait for Clk_period;
		Addr <=  "0100101000101";
		Trees_din <= x"66fff808";
		wait for Clk_period;
		Addr <=  "0100101000110";
		Trees_din <= x"adff6204";
		wait for Clk_period;
		Addr <=  "0100101000111";
		Trees_din <= x"fff32531";
		wait for Clk_period;
		Addr <=  "0100101001000";
		Trees_din <= x"00602531";
		wait for Clk_period;
		Addr <=  "0100101001001";
		Trees_din <= x"0fff2404";
		wait for Clk_period;
		Addr <=  "0100101001010";
		Trees_din <= x"00382531";
		wait for Clk_period;
		Addr <=  "0100101001011";
		Trees_din <= x"ffad2531";
		wait for Clk_period;
		Addr <=  "0100101001100";
		Trees_din <= x"bfff4030";
		wait for Clk_period;
		Addr <=  "0100101001101";
		Trees_din <= x"a9ffcb28";
		wait for Clk_period;
		Addr <=  "0100101001110";
		Trees_din <= x"8dfe9014";
		wait for Clk_period;
		Addr <=  "0100101001111";
		Trees_din <= x"b4fe850c";
		wait for Clk_period;
		Addr <=  "0100101010000";
		Trees_din <= x"cafe6008";
		wait for Clk_period;
		Addr <=  "0100101010001";
		Trees_din <= x"93ff7204";
		wait for Clk_period;
		Addr <=  "0100101010010";
		Trees_din <= x"005c2605";
		wait for Clk_period;
		Addr <=  "0100101010011";
		Trees_din <= x"ffff2605";
		wait for Clk_period;
		Addr <=  "0100101010100";
		Trees_din <= x"ffd32605";
		wait for Clk_period;
		Addr <=  "0100101010101";
		Trees_din <= x"01fef404";
		wait for Clk_period;
		Addr <=  "0100101010110";
		Trees_din <= x"ff9f2605";
		wait for Clk_period;
		Addr <=  "0100101010111";
		Trees_din <= x"00122605";
		wait for Clk_period;
		Addr <=  "0100101011000";
		Trees_din <= x"8effbb08";
		wait for Clk_period;
		Addr <=  "0100101011001";
		Trees_din <= x"dc009b04";
		wait for Clk_period;
		Addr <=  "0100101011010";
		Trees_din <= x"ffa92605";
		wait for Clk_period;
		Addr <=  "0100101011011";
		Trees_din <= x"003b2605";
		wait for Clk_period;
		Addr <=  "0100101011100";
		Trees_din <= x"abffbd04";
		wait for Clk_period;
		Addr <=  "0100101011101";
		Trees_din <= x"ffe32605";
		wait for Clk_period;
		Addr <=  "0100101011110";
		Trees_din <= x"f7ff2e04";
		wait for Clk_period;
		Addr <=  "0100101011111";
		Trees_din <= x"000c2605";
		wait for Clk_period;
		Addr <=  "0100101100000";
		Trees_din <= x"005f2605";
		wait for Clk_period;
		Addr <=  "0100101100001";
		Trees_din <= x"27000804";
		wait for Clk_period;
		Addr <=  "0100101100010";
		Trees_din <= x"ffa02605";
		wait for Clk_period;
		Addr <=  "0100101100011";
		Trees_din <= x"00152605";
		wait for Clk_period;
		Addr <=  "0100101100100";
		Trees_din <= x"c5ff3120";
		wait for Clk_period;
		Addr <=  "0100101100101";
		Trees_din <= x"28ff310c";
		wait for Clk_period;
		Addr <=  "0100101100110";
		Trees_din <= x"1afe2904";
		wait for Clk_period;
		Addr <=  "0100101100111";
		Trees_din <= x"00302605";
		wait for Clk_period;
		Addr <=  "0100101101000";
		Trees_din <= x"b5ff3104";
		wait for Clk_period;
		Addr <=  "0100101101001";
		Trees_din <= x"ff8c2605";
		wait for Clk_period;
		Addr <=  "0100101101010";
		Trees_din <= x"ffe92605";
		wait for Clk_period;
		Addr <=  "0100101101011";
		Trees_din <= x"71ff3d0c";
		wait for Clk_period;
		Addr <=  "0100101101100";
		Trees_din <= x"7efec004";
		wait for Clk_period;
		Addr <=  "0100101101101";
		Trees_din <= x"fff82605";
		wait for Clk_period;
		Addr <=  "0100101101110";
		Trees_din <= x"86feee04";
		wait for Clk_period;
		Addr <=  "0100101101111";
		Trees_din <= x"00142605";
		wait for Clk_period;
		Addr <=  "0100101110000";
		Trees_din <= x"00752605";
		wait for Clk_period;
		Addr <=  "0100101110001";
		Trees_din <= x"28ff5104";
		wait for Clk_period;
		Addr <=  "0100101110010";
		Trees_din <= x"00392605";
		wait for Clk_period;
		Addr <=  "0100101110011";
		Trees_din <= x"ffb12605";
		wait for Clk_period;
		Addr <=  "0100101110100";
		Trees_din <= x"0a007a08";
		wait for Clk_period;
		Addr <=  "0100101110101";
		Trees_din <= x"4ffed804";
		wait for Clk_period;
		Addr <=  "0100101110110";
		Trees_din <= x"ffed2605";
		wait for Clk_period;
		Addr <=  "0100101110111";
		Trees_din <= x"ff812605";
		wait for Clk_period;
		Addr <=  "0100101111000";
		Trees_din <= x"39ff7708";
		wait for Clk_period;
		Addr <=  "0100101111001";
		Trees_din <= x"43ff9204";
		wait for Clk_period;
		Addr <=  "0100101111010";
		Trees_din <= x"ffe22605";
		wait for Clk_period;
		Addr <=  "0100101111011";
		Trees_din <= x"004e2605";
		wait for Clk_period;
		Addr <=  "0100101111100";
		Trees_din <= x"00002a08";
		wait for Clk_period;
		Addr <=  "0100101111101";
		Trees_din <= x"8a004704";
		wait for Clk_period;
		Addr <=  "0100101111110";
		Trees_din <= x"ff962605";
		wait for Clk_period;
		Addr <=  "0100101111111";
		Trees_din <= x"ffe62605";
		wait for Clk_period;
		Addr <=  "0100110000000";
		Trees_din <= x"00142605";
		wait for Clk_period;
		Addr <=  "0100110000001";
		Trees_din <= x"0fff3124";
		wait for Clk_period;
		Addr <=  "0100110000010";
		Trees_din <= x"f7ff2e0c";
		wait for Clk_period;
		Addr <=  "0100110000011";
		Trees_din <= x"dc00b708";
		wait for Clk_period;
		Addr <=  "0100110000100";
		Trees_din <= x"27005104";
		wait for Clk_period;
		Addr <=  "0100110000101";
		Trees_din <= x"ff9a26c9";
		wait for Clk_period;
		Addr <=  "0100110000110";
		Trees_din <= x"000c26c9";
		wait for Clk_period;
		Addr <=  "0100110000111";
		Trees_din <= x"003b26c9";
		wait for Clk_period;
		Addr <=  "0100110001000";
		Trees_din <= x"25ffb404";
		wait for Clk_period;
		Addr <=  "0100110001001";
		Trees_din <= x"ffdc26c9";
		wait for Clk_period;
		Addr <=  "0100110001010";
		Trees_din <= x"67ffba10";
		wait for Clk_period;
		Addr <=  "0100110001011";
		Trees_din <= x"71ff7a08";
		wait for Clk_period;
		Addr <=  "0100110001100";
		Trees_din <= x"ec001d04";
		wait for Clk_period;
		Addr <=  "0100110001101";
		Trees_din <= x"006a26c9";
		wait for Clk_period;
		Addr <=  "0100110001110";
		Trees_din <= x"000f26c9";
		wait for Clk_period;
		Addr <=  "0100110001111";
		Trees_din <= x"42ffa804";
		wait for Clk_period;
		Addr <=  "0100110010000";
		Trees_din <= x"ffbe26c9";
		wait for Clk_period;
		Addr <=  "0100110010001";
		Trees_din <= x"003926c9";
		wait for Clk_period;
		Addr <=  "0100110010010";
		Trees_din <= x"ffe026c9";
		wait for Clk_period;
		Addr <=  "0100110010011";
		Trees_din <= x"30ffb50c";
		wait for Clk_period;
		Addr <=  "0100110010100";
		Trees_din <= x"95ffa708";
		wait for Clk_period;
		Addr <=  "0100110010101";
		Trees_din <= x"7fffce04";
		wait for Clk_period;
		Addr <=  "0100110010110";
		Trees_din <= x"ff7f26c9";
		wait for Clk_period;
		Addr <=  "0100110010111";
		Trees_din <= x"fffe26c9";
		wait for Clk_period;
		Addr <=  "0100110011000";
		Trees_din <= x"001326c9";
		wait for Clk_period;
		Addr <=  "0100110011001";
		Trees_din <= x"ac003718";
		wait for Clk_period;
		Addr <=  "0100110011010";
		Trees_din <= x"5a001a0c";
		wait for Clk_period;
		Addr <=  "0100110011011";
		Trees_din <= x"5bff5004";
		wait for Clk_period;
		Addr <=  "0100110011100";
		Trees_din <= x"ffc426c9";
		wait for Clk_period;
		Addr <=  "0100110011101";
		Trees_din <= x"4cff4a04";
		wait for Clk_period;
		Addr <=  "0100110011110";
		Trees_din <= x"fff926c9";
		wait for Clk_period;
		Addr <=  "0100110011111";
		Trees_din <= x"005326c9";
		wait for Clk_period;
		Addr <=  "0100110100000";
		Trees_din <= x"19ffad08";
		wait for Clk_period;
		Addr <=  "0100110100001";
		Trees_din <= x"dc00be04";
		wait for Clk_period;
		Addr <=  "0100110100010";
		Trees_din <= x"ff8d26c9";
		wait for Clk_period;
		Addr <=  "0100110100011";
		Trees_din <= x"001426c9";
		wait for Clk_period;
		Addr <=  "0100110100100";
		Trees_din <= x"001426c9";
		wait for Clk_period;
		Addr <=  "0100110100101";
		Trees_din <= x"ac005c0c";
		wait for Clk_period;
		Addr <=  "0100110100110";
		Trees_din <= x"a9ffac08";
		wait for Clk_period;
		Addr <=  "0100110100111";
		Trees_din <= x"be000c04";
		wait for Clk_period;
		Addr <=  "0100110101000";
		Trees_din <= x"006b26c9";
		wait for Clk_period;
		Addr <=  "0100110101001";
		Trees_din <= x"000426c9";
		wait for Clk_period;
		Addr <=  "0100110101010";
		Trees_din <= x"ffe826c9";
		wait for Clk_period;
		Addr <=  "0100110101011";
		Trees_din <= x"faff7f08";
		wait for Clk_period;
		Addr <=  "0100110101100";
		Trees_din <= x"e4fe2c04";
		wait for Clk_period;
		Addr <=  "0100110101101";
		Trees_din <= x"002826c9";
		wait for Clk_period;
		Addr <=  "0100110101110";
		Trees_din <= x"ffa426c9";
		wait for Clk_period;
		Addr <=  "0100110101111";
		Trees_din <= x"39ffa404";
		wait for Clk_period;
		Addr <=  "0100110110000";
		Trees_din <= x"004326c9";
		wait for Clk_period;
		Addr <=  "0100110110001";
		Trees_din <= x"ffd626c9";
		wait for Clk_period;
		Addr <=  "0100110110010";
		Trees_din <= x"aaff7330";
		wait for Clk_period;
		Addr <=  "0100110110011";
		Trees_din <= x"b4fe9a18";
		wait for Clk_period;
		Addr <=  "0100110110100";
		Trees_din <= x"09fff210";
		wait for Clk_period;
		Addr <=  "0100110110101";
		Trees_din <= x"60ffbc0c";
		wait for Clk_period;
		Addr <=  "0100110110110";
		Trees_din <= x"4cff0704";
		wait for Clk_period;
		Addr <=  "0100110110111";
		Trees_din <= x"fff6279d";
		wait for Clk_period;
		Addr <=  "0100110111000";
		Trees_din <= x"c8000a04";
		wait for Clk_period;
		Addr <=  "0100110111001";
		Trees_din <= x"0015279d";
		wait for Clk_period;
		Addr <=  "0100110111010";
		Trees_din <= x"0064279d";
		wait for Clk_period;
		Addr <=  "0100110111011";
		Trees_din <= x"ffe0279d";
		wait for Clk_period;
		Addr <=  "0100110111100";
		Trees_din <= x"87ff7304";
		wait for Clk_period;
		Addr <=  "0100110111101";
		Trees_din <= x"ffb1279d";
		wait for Clk_period;
		Addr <=  "0100110111110";
		Trees_din <= x"0024279d";
		wait for Clk_period;
		Addr <=  "0100110111111";
		Trees_din <= x"0cfe2e0c";
		wait for Clk_period;
		Addr <=  "0100111000000";
		Trees_din <= x"daffbc04";
		wait for Clk_period;
		Addr <=  "0100111000001";
		Trees_din <= x"ffbc279d";
		wait for Clk_period;
		Addr <=  "0100111000010";
		Trees_din <= x"afffd704";
		wait for Clk_period;
		Addr <=  "0100111000011";
		Trees_din <= x"fff1279d";
		wait for Clk_period;
		Addr <=  "0100111000100";
		Trees_din <= x"0047279d";
		wait for Clk_period;
		Addr <=  "0100111000101";
		Trees_din <= x"e7feff04";
		wait for Clk_period;
		Addr <=  "0100111000110";
		Trees_din <= x"0000279d";
		wait for Clk_period;
		Addr <=  "0100111000111";
		Trees_din <= x"a6fee404";
		wait for Clk_period;
		Addr <=  "0100111001000";
		Trees_din <= x"fff3279d";
		wait for Clk_period;
		Addr <=  "0100111001001";
		Trees_din <= x"ff85279d";
		wait for Clk_period;
		Addr <=  "0100111001010";
		Trees_din <= x"e2ff231c";
		wait for Clk_period;
		Addr <=  "0100111001011";
		Trees_din <= x"0fffaa10";
		wait for Clk_period;
		Addr <=  "0100111001100";
		Trees_din <= x"2cff3904";
		wait for Clk_period;
		Addr <=  "0100111001101";
		Trees_din <= x"ffda279d";
		wait for Clk_period;
		Addr <=  "0100111001110";
		Trees_din <= x"de006208";
		wait for Clk_period;
		Addr <=  "0100111001111";
		Trees_din <= x"aefe9404";
		wait for Clk_period;
		Addr <=  "0100111010000";
		Trees_din <= x"000d279d";
		wait for Clk_period;
		Addr <=  "0100111010001";
		Trees_din <= x"0063279d";
		wait for Clk_period;
		Addr <=  "0100111010010";
		Trees_din <= x"fff0279d";
		wait for Clk_period;
		Addr <=  "0100111010011";
		Trees_din <= x"de008808";
		wait for Clk_period;
		Addr <=  "0100111010100";
		Trees_din <= x"e8ff4c04";
		wait for Clk_period;
		Addr <=  "0100111010101";
		Trees_din <= x"0015279d";
		wait for Clk_period;
		Addr <=  "0100111010110";
		Trees_din <= x"ffa4279d";
		wait for Clk_period;
		Addr <=  "0100111010111";
		Trees_din <= x"003a279d";
		wait for Clk_period;
		Addr <=  "0100111011000";
		Trees_din <= x"e8ff9614";
		wait for Clk_period;
		Addr <=  "0100111011001";
		Trees_din <= x"01fea408";
		wait for Clk_period;
		Addr <=  "0100111011010";
		Trees_din <= x"a7ffab04";
		wait for Clk_period;
		Addr <=  "0100111011011";
		Trees_din <= x"ffb1279d";
		wait for Clk_period;
		Addr <=  "0100111011100";
		Trees_din <= x"fffe279d";
		wait for Clk_period;
		Addr <=  "0100111011101";
		Trees_din <= x"1eff9c04";
		wait for Clk_period;
		Addr <=  "0100111011110";
		Trees_din <= x"ffda279d";
		wait for Clk_period;
		Addr <=  "0100111011111";
		Trees_din <= x"2affc504";
		wait for Clk_period;
		Addr <=  "0100111100000";
		Trees_din <= x"0006279d";
		wait for Clk_period;
		Addr <=  "0100111100001";
		Trees_din <= x"005e279d";
		wait for Clk_period;
		Addr <=  "0100111100010";
		Trees_din <= x"0eff5308";
		wait for Clk_period;
		Addr <=  "0100111100011";
		Trees_din <= x"e4fe6904";
		wait for Clk_period;
		Addr <=  "0100111100100";
		Trees_din <= x"ffea279d";
		wait for Clk_period;
		Addr <=  "0100111100101";
		Trees_din <= x"ff90279d";
		wait for Clk_period;
		Addr <=  "0100111100110";
		Trees_din <= x"0014279d";
		wait for Clk_period;
		Addr <=  "0100111100111";
		Trees_din <= x"bfff4030";
		wait for Clk_period;
		Addr <=  "0100111101000";
		Trees_din <= x"0dff7e1c";
		wait for Clk_period;
		Addr <=  "0100111101001";
		Trees_din <= x"3cfed508";
		wait for Clk_period;
		Addr <=  "0100111101010";
		Trees_din <= x"bdff6604";
		wait for Clk_period;
		Addr <=  "0100111101011";
		Trees_din <= x"00222859";
		wait for Clk_period;
		Addr <=  "0100111101100";
		Trees_din <= x"ffad2859";
		wait for Clk_period;
		Addr <=  "0100111101101";
		Trees_din <= x"a9ffcb0c";
		wait for Clk_period;
		Addr <=  "0100111101110";
		Trees_din <= x"4bff4d08";
		wait for Clk_period;
		Addr <=  "0100111101111";
		Trees_din <= x"36ffc004";
		wait for Clk_period;
		Addr <=  "0100111110000";
		Trees_din <= x"00592859";
		wait for Clk_period;
		Addr <=  "0100111110001";
		Trees_din <= x"ffed2859";
		wait for Clk_period;
		Addr <=  "0100111110010";
		Trees_din <= x"ffec2859";
		wait for Clk_period;
		Addr <=  "0100111110011";
		Trees_din <= x"e3fecd04";
		wait for Clk_period;
		Addr <=  "0100111110100";
		Trees_din <= x"ffc02859";
		wait for Clk_period;
		Addr <=  "0100111110101";
		Trees_din <= x"00122859";
		wait for Clk_period;
		Addr <=  "0100111110110";
		Trees_din <= x"04007908";
		wait for Clk_period;
		Addr <=  "0100111110111";
		Trees_din <= x"c5ff2404";
		wait for Clk_period;
		Addr <=  "0100111111000";
		Trees_din <= x"00002859";
		wait for Clk_period;
		Addr <=  "0100111111001";
		Trees_din <= x"ff972859";
		wait for Clk_period;
		Addr <=  "0100111111010";
		Trees_din <= x"88ffee04";
		wait for Clk_period;
		Addr <=  "0100111111011";
		Trees_din <= x"ffd12859";
		wait for Clk_period;
		Addr <=  "0100111111100";
		Trees_din <= x"97feb504";
		wait for Clk_period;
		Addr <=  "0100111111101";
		Trees_din <= x"00512859";
		wait for Clk_period;
		Addr <=  "0100111111110";
		Trees_din <= x"00032859";
		wait for Clk_period;
		Addr <=  "0100111111111";
		Trees_din <= x"c5ff3118";
		wait for Clk_period;
		Addr <=  "0101000000000";
		Trees_din <= x"28ff3108";
		wait for Clk_period;
		Addr <=  "0101000000001";
		Trees_din <= x"59feec04";
		wait for Clk_period;
		Addr <=  "0101000000010";
		Trees_din <= x"00212859";
		wait for Clk_period;
		Addr <=  "0101000000011";
		Trees_din <= x"ff9d2859";
		wait for Clk_period;
		Addr <=  "0101000000100";
		Trees_din <= x"2aff8704";
		wait for Clk_period;
		Addr <=  "0101000000101";
		Trees_din <= x"ffd72859";
		wait for Clk_period;
		Addr <=  "0101000000110";
		Trees_din <= x"f1ffc508";
		wait for Clk_period;
		Addr <=  "0101000000111";
		Trees_din <= x"c9fff704";
		wait for Clk_period;
		Addr <=  "0101000001000";
		Trees_din <= x"005c2859";
		wait for Clk_period;
		Addr <=  "0101000001001";
		Trees_din <= x"fffa2859";
		wait for Clk_period;
		Addr <=  "0101000001010";
		Trees_din <= x"ffed2859";
		wait for Clk_period;
		Addr <=  "0101000001011";
		Trees_din <= x"8a00350c";
		wait for Clk_period;
		Addr <=  "0101000001100";
		Trees_din <= x"ce001e08";
		wait for Clk_period;
		Addr <=  "0101000001101";
		Trees_din <= x"3eff2c04";
		wait for Clk_period;
		Addr <=  "0101000001110";
		Trees_din <= x"ffd92859";
		wait for Clk_period;
		Addr <=  "0101000001111";
		Trees_din <= x"ff7f2859";
		wait for Clk_period;
		Addr <=  "0101000010000";
		Trees_din <= x"001a2859";
		wait for Clk_period;
		Addr <=  "0101000010001";
		Trees_din <= x"81ff7108";
		wait for Clk_period;
		Addr <=  "0101000010010";
		Trees_din <= x"a1ff6904";
		wait for Clk_period;
		Addr <=  "0101000010011";
		Trees_din <= x"fffb2859";
		wait for Clk_period;
		Addr <=  "0101000010100";
		Trees_din <= x"00452859";
		wait for Clk_period;
		Addr <=  "0101000010101";
		Trees_din <= x"ffc82859";
		wait for Clk_period;
		Addr <=  "0101000010110";
		Trees_din <= x"2cff6a18";
		wait for Clk_period;
		Addr <=  "0101000010111";
		Trees_din <= x"3000110c";
		wait for Clk_period;
		Addr <=  "0101000011000";
		Trees_din <= x"97fe7004";
		wait for Clk_period;
		Addr <=  "0101000011001";
		Trees_din <= x"001228fd";
		wait for Clk_period;
		Addr <=  "0101000011010";
		Trees_din <= x"dc006204";
		wait for Clk_period;
		Addr <=  "0101000011011";
		Trees_din <= x"ff8b28fd";
		wait for Clk_period;
		Addr <=  "0101000011100";
		Trees_din <= x"fff328fd";
		wait for Clk_period;
		Addr <=  "0101000011101";
		Trees_din <= x"08004a04";
		wait for Clk_period;
		Addr <=  "0101000011110";
		Trees_din <= x"ffc328fd";
		wait for Clk_period;
		Addr <=  "0101000011111";
		Trees_din <= x"f0ff0c04";
		wait for Clk_period;
		Addr <=  "0101000100000";
		Trees_din <= x"004128fd";
		wait for Clk_period;
		Addr <=  "0101000100001";
		Trees_din <= x"ffed28fd";
		wait for Clk_period;
		Addr <=  "0101000100010";
		Trees_din <= x"88ffd010";
		wait for Clk_period;
		Addr <=  "0101000100011";
		Trees_din <= x"c7fea508";
		wait for Clk_period;
		Addr <=  "0101000100100";
		Trees_din <= x"f3fefd04";
		wait for Clk_period;
		Addr <=  "0101000100101";
		Trees_din <= x"ffe628fd";
		wait for Clk_period;
		Addr <=  "0101000100110";
		Trees_din <= x"003928fd";
		wait for Clk_period;
		Addr <=  "0101000100111";
		Trees_din <= x"8dff3504";
		wait for Clk_period;
		Addr <=  "0101000101000";
		Trees_din <= x"ff9328fd";
		wait for Clk_period;
		Addr <=  "0101000101001";
		Trees_din <= x"ffe728fd";
		wait for Clk_period;
		Addr <=  "0101000101010";
		Trees_din <= x"71ff3d10";
		wait for Clk_period;
		Addr <=  "0101000101011";
		Trees_din <= x"8c007c0c";
		wait for Clk_period;
		Addr <=  "0101000101100";
		Trees_din <= x"2b005708";
		wait for Clk_period;
		Addr <=  "0101000101101";
		Trees_din <= x"36ff8604";
		wait for Clk_period;
		Addr <=  "0101000101110";
		Trees_din <= x"005128fd";
		wait for Clk_period;
		Addr <=  "0101000101111";
		Trees_din <= x"000828fd";
		wait for Clk_period;
		Addr <=  "0101000110000";
		Trees_din <= x"ffd728fd";
		wait for Clk_period;
		Addr <=  "0101000110001";
		Trees_din <= x"ffdf28fd";
		wait for Clk_period;
		Addr <=  "0101000110010";
		Trees_din <= x"fb001d10";
		wait for Clk_period;
		Addr <=  "0101000110011";
		Trees_din <= x"60ff2908";
		wait for Clk_period;
		Addr <=  "0101000110100";
		Trees_din <= x"ac003104";
		wait for Clk_period;
		Addr <=  "0101000110101";
		Trees_din <= x"fff328fd";
		wait for Clk_period;
		Addr <=  "0101000110110";
		Trees_din <= x"004428fd";
		wait for Clk_period;
		Addr <=  "0101000110111";
		Trees_din <= x"2a00fe04";
		wait for Clk_period;
		Addr <=  "0101000111000";
		Trees_din <= x"ffa428fd";
		wait for Clk_period;
		Addr <=  "0101000111001";
		Trees_din <= x"001328fd";
		wait for Clk_period;
		Addr <=  "0101000111010";
		Trees_din <= x"c1fea604";
		wait for Clk_period;
		Addr <=  "0101000111011";
		Trees_din <= x"fff328fd";
		wait for Clk_period;
		Addr <=  "0101000111100";
		Trees_din <= x"92ff1f04";
		wait for Clk_period;
		Addr <=  "0101000111101";
		Trees_din <= x"001728fd";
		wait for Clk_period;
		Addr <=  "0101000111110";
		Trees_din <= x"005e28fd";
		wait for Clk_period;
		Addr <=  "0101000111111";
		Trees_din <= x"9cff7c2c";
		wait for Clk_period;
		Addr <=  "0101001000000";
		Trees_din <= x"faff7a10";
		wait for Clk_period;
		Addr <=  "0101001000001";
		Trees_din <= x"59feb504";
		wait for Clk_period;
		Addr <=  "0101001000010";
		Trees_din <= x"002429d1";
		wait for Clk_period;
		Addr <=  "0101001000011";
		Trees_din <= x"6bfe3104";
		wait for Clk_period;
		Addr <=  "0101001000100";
		Trees_din <= x"000629d1";
		wait for Clk_period;
		Addr <=  "0101001000101";
		Trees_din <= x"0a00b904";
		wait for Clk_period;
		Addr <=  "0101001000110";
		Trees_din <= x"ff8329d1";
		wait for Clk_period;
		Addr <=  "0101001000111";
		Trees_din <= x"ffde29d1";
		wait for Clk_period;
		Addr <=  "0101001001000";
		Trees_din <= x"efffa014";
		wait for Clk_period;
		Addr <=  "0101001001001";
		Trees_din <= x"00ff7208";
		wait for Clk_period;
		Addr <=  "0101001001010";
		Trees_din <= x"11ff7804";
		wait for Clk_period;
		Addr <=  "0101001001011";
		Trees_din <= x"ffb829d1";
		wait for Clk_period;
		Addr <=  "0101001001100";
		Trees_din <= x"001d29d1";
		wait for Clk_period;
		Addr <=  "0101001001101";
		Trees_din <= x"64ff2a08";
		wait for Clk_period;
		Addr <=  "0101001001110";
		Trees_din <= x"0efed004";
		wait for Clk_period;
		Addr <=  "0101001001111";
		Trees_din <= x"000729d1";
		wait for Clk_period;
		Addr <=  "0101001010000";
		Trees_din <= x"006429d1";
		wait for Clk_period;
		Addr <=  "0101001010001";
		Trees_din <= x"fff929d1";
		wait for Clk_period;
		Addr <=  "0101001010010";
		Trees_din <= x"ccff6004";
		wait for Clk_period;
		Addr <=  "0101001010011";
		Trees_din <= x"000329d1";
		wait for Clk_period;
		Addr <=  "0101001010100";
		Trees_din <= x"ffa629d1";
		wait for Clk_period;
		Addr <=  "0101001010101";
		Trees_din <= x"28ff291c";
		wait for Clk_period;
		Addr <=  "0101001010110";
		Trees_din <= x"bffeeb0c";
		wait for Clk_period;
		Addr <=  "0101001010111";
		Trees_din <= x"35fefb08";
		wait for Clk_period;
		Addr <=  "0101001011000";
		Trees_din <= x"0efeba04";
		wait for Clk_period;
		Addr <=  "0101001011001";
		Trees_din <= x"000329d1";
		wait for Clk_period;
		Addr <=  "0101001011010";
		Trees_din <= x"005229d1";
		wait for Clk_period;
		Addr <=  "0101001011011";
		Trees_din <= x"ffd329d1";
		wait for Clk_period;
		Addr <=  "0101001011100";
		Trees_din <= x"01fe3a08";
		wait for Clk_period;
		Addr <=  "0101001011101";
		Trees_din <= x"1cff3004";
		wait for Clk_period;
		Addr <=  "0101001011110";
		Trees_din <= x"002f29d1";
		wait for Clk_period;
		Addr <=  "0101001011111";
		Trees_din <= x"ffe929d1";
		wait for Clk_period;
		Addr <=  "0101001100000";
		Trees_din <= x"42ffe204";
		wait for Clk_period;
		Addr <=  "0101001100001";
		Trees_din <= x"ff9629d1";
		wait for Clk_period;
		Addr <=  "0101001100010";
		Trees_din <= x"fff929d1";
		wait for Clk_period;
		Addr <=  "0101001100011";
		Trees_din <= x"d3fef014";
		wait for Clk_period;
		Addr <=  "0101001100100";
		Trees_din <= x"a3ff7608";
		wait for Clk_period;
		Addr <=  "0101001100101";
		Trees_din <= x"82ff7104";
		wait for Clk_period;
		Addr <=  "0101001100110";
		Trees_din <= x"ffa929d1";
		wait for Clk_period;
		Addr <=  "0101001100111";
		Trees_din <= x"001129d1";
		wait for Clk_period;
		Addr <=  "0101001101000";
		Trees_din <= x"80ff8304";
		wait for Clk_period;
		Addr <=  "0101001101001";
		Trees_din <= x"ffe229d1";
		wait for Clk_period;
		Addr <=  "0101001101010";
		Trees_din <= x"12ffbd04";
		wait for Clk_period;
		Addr <=  "0101001101011";
		Trees_din <= x"fffa29d1";
		wait for Clk_period;
		Addr <=  "0101001101100";
		Trees_din <= x"005429d1";
		wait for Clk_period;
		Addr <=  "0101001101101";
		Trees_din <= x"4bff3b0c";
		wait for Clk_period;
		Addr <=  "0101001101110";
		Trees_din <= x"2cff7304";
		wait for Clk_period;
		Addr <=  "0101001101111";
		Trees_din <= x"fffa29d1";
		wait for Clk_period;
		Addr <=  "0101001110000";
		Trees_din <= x"7bff9b04";
		wait for Clk_period;
		Addr <=  "0101001110001";
		Trees_din <= x"005f29d1";
		wait for Clk_period;
		Addr <=  "0101001110010";
		Trees_din <= x"000129d1";
		wait for Clk_period;
		Addr <=  "0101001110011";
		Trees_din <= x"ffee29d1";
		wait for Clk_period;
		Addr <=  "0101001110100";
		Trees_din <= x"64fede20";
		wait for Clk_period;
		Addr <=  "0101001110101";
		Trees_din <= x"de00621c";
		wait for Clk_period;
		Addr <=  "0101001110110";
		Trees_din <= x"c1febc10";
		wait for Clk_period;
		Addr <=  "0101001110111";
		Trees_din <= x"1b004f0c";
		wait for Clk_period;
		Addr <=  "0101001111000";
		Trees_din <= x"f3ff5f08";
		wait for Clk_period;
		Addr <=  "0101001111001";
		Trees_din <= x"a0ff4404";
		wait for Clk_period;
		Addr <=  "0101001111010";
		Trees_din <= x"ffad2a85";
		wait for Clk_period;
		Addr <=  "0101001111011";
		Trees_din <= x"fff32a85";
		wait for Clk_period;
		Addr <=  "0101001111100";
		Trees_din <= x"00132a85";
		wait for Clk_period;
		Addr <=  "0101001111101";
		Trees_din <= x"00412a85";
		wait for Clk_period;
		Addr <=  "0101001111110";
		Trees_din <= x"67ff8508";
		wait for Clk_period;
		Addr <=  "0101001111111";
		Trees_din <= x"31003804";
		wait for Clk_period;
		Addr <=  "0101010000000";
		Trees_din <= x"00662a85";
		wait for Clk_period;
		Addr <=  "0101010000001";
		Trees_din <= x"00062a85";
		wait for Clk_period;
		Addr <=  "0101010000010";
		Trees_din <= x"fff82a85";
		wait for Clk_period;
		Addr <=  "0101010000011";
		Trees_din <= x"ffc72a85";
		wait for Clk_period;
		Addr <=  "0101010000100";
		Trees_din <= x"c5ff2d1c";
		wait for Clk_period;
		Addr <=  "0101010000101";
		Trees_din <= x"f7ff2e0c";
		wait for Clk_period;
		Addr <=  "0101010000110";
		Trees_din <= x"11ffc908";
		wait for Clk_period;
		Addr <=  "0101010000111";
		Trees_din <= x"12ff8e04";
		wait for Clk_period;
		Addr <=  "0101010001000";
		Trees_din <= x"fff92a85";
		wait for Clk_period;
		Addr <=  "0101010001001";
		Trees_din <= x"ff9a2a85";
		wait for Clk_period;
		Addr <=  "0101010001010";
		Trees_din <= x"001e2a85";
		wait for Clk_period;
		Addr <=  "0101010001011";
		Trees_din <= x"8effcb04";
		wait for Clk_period;
		Addr <=  "0101010001100";
		Trees_din <= x"ffd52a85";
		wait for Clk_period;
		Addr <=  "0101010001101";
		Trees_din <= x"f3febe04";
		wait for Clk_period;
		Addr <=  "0101010001110";
		Trees_din <= x"fff22a85";
		wait for Clk_period;
		Addr <=  "0101010001111";
		Trees_din <= x"1f006f04";
		wait for Clk_period;
		Addr <=  "0101010010000";
		Trees_din <= x"005d2a85";
		wait for Clk_period;
		Addr <=  "0101010010001";
		Trees_din <= x"fff92a85";
		wait for Clk_period;
		Addr <=  "0101010010010";
		Trees_din <= x"83fe9208";
		wait for Clk_period;
		Addr <=  "0101010010011";
		Trees_din <= x"dcff5604";
		wait for Clk_period;
		Addr <=  "0101010010100";
		Trees_din <= x"003f2a85";
		wait for Clk_period;
		Addr <=  "0101010010101";
		Trees_din <= x"fff52a85";
		wait for Clk_period;
		Addr <=  "0101010010110";
		Trees_din <= x"1cfee608";
		wait for Clk_period;
		Addr <=  "0101010010111";
		Trees_din <= x"a2ff9004";
		wait for Clk_period;
		Addr <=  "0101010011000";
		Trees_din <= x"00392a85";
		wait for Clk_period;
		Addr <=  "0101010011001";
		Trees_din <= x"ffda2a85";
		wait for Clk_period;
		Addr <=  "0101010011010";
		Trees_din <= x"b7ff1b08";
		wait for Clk_period;
		Addr <=  "0101010011011";
		Trees_din <= x"ebff0504";
		wait for Clk_period;
		Addr <=  "0101010011100";
		Trees_din <= x"ffde2a85";
		wait for Clk_period;
		Addr <=  "0101010011101";
		Trees_din <= x"00202a85";
		wait for Clk_period;
		Addr <=  "0101010011110";
		Trees_din <= x"4cffe504";
		wait for Clk_period;
		Addr <=  "0101010011111";
		Trees_din <= x"ff902a85";
		wait for Clk_period;
		Addr <=  "0101010100000";
		Trees_din <= x"fff92a85";
		wait for Clk_period;
		Addr <=  "0101010100001";
		Trees_din <= x"8dfe9024";
		wait for Clk_period;
		Addr <=  "0101010100010";
		Trees_din <= x"89015520";
		wait for Clk_period;
		Addr <=  "0101010100011";
		Trees_din <= x"32fe4608";
		wait for Clk_period;
		Addr <=  "0101010100100";
		Trees_din <= x"53ffb604";
		wait for Clk_period;
		Addr <=  "0101010100101";
		Trees_din <= x"ffeb2b39";
		wait for Clk_period;
		Addr <=  "0101010100110";
		Trees_din <= x"00392b39";
		wait for Clk_period;
		Addr <=  "0101010100111";
		Trees_din <= x"28ff5a0c";
		wait for Clk_period;
		Addr <=  "0101010101000";
		Trees_din <= x"89005d04";
		wait for Clk_period;
		Addr <=  "0101010101001";
		Trees_din <= x"ff8a2b39";
		wait for Clk_period;
		Addr <=  "0101010101010";
		Trees_din <= x"34000904";
		wait for Clk_period;
		Addr <=  "0101010101011";
		Trees_din <= x"00102b39";
		wait for Clk_period;
		Addr <=  "0101010101100";
		Trees_din <= x"ffbb2b39";
		wait for Clk_period;
		Addr <=  "0101010101101";
		Trees_din <= x"4fffb308";
		wait for Clk_period;
		Addr <=  "0101010101110";
		Trees_din <= x"faff9f04";
		wait for Clk_period;
		Addr <=  "0101010101111";
		Trees_din <= x"ffab2b39";
		wait for Clk_period;
		Addr <=  "0101010110000";
		Trees_din <= x"000b2b39";
		wait for Clk_period;
		Addr <=  "0101010110001";
		Trees_din <= x"00262b39";
		wait for Clk_period;
		Addr <=  "0101010110010";
		Trees_din <= x"00352b39";
		wait for Clk_period;
		Addr <=  "0101010110011";
		Trees_din <= x"97fee518";
		wait for Clk_period;
		Addr <=  "0101010110100";
		Trees_din <= x"66ffaf08";
		wait for Clk_period;
		Addr <=  "0101010110101";
		Trees_din <= x"57feb704";
		wait for Clk_period;
		Addr <=  "0101010110110";
		Trees_din <= x"001e2b39";
		wait for Clk_period;
		Addr <=  "0101010110111";
		Trees_din <= x"ffbf2b39";
		wait for Clk_period;
		Addr <=  "0101010111000";
		Trees_din <= x"45ff3d0c";
		wait for Clk_period;
		Addr <=  "0101010111001";
		Trees_din <= x"8effc904";
		wait for Clk_period;
		Addr <=  "0101010111010";
		Trees_din <= x"fffe2b39";
		wait for Clk_period;
		Addr <=  "0101010111011";
		Trees_din <= x"7aff4d04";
		wait for Clk_period;
		Addr <=  "0101010111100";
		Trees_din <= x"00142b39";
		wait for Clk_period;
		Addr <=  "0101010111101";
		Trees_din <= x"00672b39";
		wait for Clk_period;
		Addr <=  "0101010111110";
		Trees_din <= x"ffee2b39";
		wait for Clk_period;
		Addr <=  "0101010111111";
		Trees_din <= x"0a00370c";
		wait for Clk_period;
		Addr <=  "0101011000000";
		Trees_din <= x"87ffbf08";
		wait for Clk_period;
		Addr <=  "0101011000001";
		Trees_din <= x"7cffdc04";
		wait for Clk_period;
		Addr <=  "0101011000010";
		Trees_din <= x"ff932b39";
		wait for Clk_period;
		Addr <=  "0101011000011";
		Trees_din <= x"ffef2b39";
		wait for Clk_period;
		Addr <=  "0101011000100";
		Trees_din <= x"00292b39";
		wait for Clk_period;
		Addr <=  "0101011000101";
		Trees_din <= x"37ff7e0c";
		wait for Clk_period;
		Addr <=  "0101011000110";
		Trees_din <= x"a9ffcb08";
		wait for Clk_period;
		Addr <=  "0101011000111";
		Trees_din <= x"85ffc004";
		wait for Clk_period;
		Addr <=  "0101011001000";
		Trees_din <= x"00022b39";
		wait for Clk_period;
		Addr <=  "0101011001001";
		Trees_din <= x"004d2b39";
		wait for Clk_period;
		Addr <=  "0101011001010";
		Trees_din <= x"ffdd2b39";
		wait for Clk_period;
		Addr <=  "0101011001011";
		Trees_din <= x"39ff8904";
		wait for Clk_period;
		Addr <=  "0101011001100";
		Trees_din <= x"00122b39";
		wait for Clk_period;
		Addr <=  "0101011001101";
		Trees_din <= x"ffb62b39";
		wait for Clk_period;
		Addr <=  "0101011001110";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  5
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"f5ff7134";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"d0009014";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"efffbb08";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"f9000d04";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"ff5700ed";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"003700ed";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"03001908";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"10002b04";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"ff7400ed";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"003700ed";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"017b00ed";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"43fef00c";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"0affbf04";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"ff9c00ed";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"1afe7f04";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"003700ed";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"036400ed";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"cdff6908";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"22005a04";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"ff9600ed";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"026e00ed";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"2cff7008";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"09fff904";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"ff8800ed";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"01ef00ed";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"ff5f00ed";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"27000524";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"82006b18";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"4afe2a08";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"17002b04";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"ff7900ed";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"015c00ed";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"5c01bf08";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"ef001704";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"ff5800ed";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"ff9b00ed";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"0800c904";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"ffa400ed";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"00ca00ed";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"ac002704";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"017b00ed";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"05005704";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"ff7100ed";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"003700ed";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"a1fdc208";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"17ff9e04";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"ff7700ed";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"01bf00ed";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"05012410";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"42feb308";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"edff5004";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"011400ed";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"ff7b00ed";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"09fdbc04";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"007000ed";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"ff6e00ed";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"9cffae04";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"ff7700ed";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"01bf00ed";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"f5ff7124";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"42ff891c";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"a7ffb818";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"e6ffe010";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"3dffbb08";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"a5feff04";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"00d401e1";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"ff8101e1";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"07ffd904";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"ff9b01e1";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"01d501e1";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"f7fec404";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"00b001e1";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"ff6d01e1";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"ff6301e1";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"4affba04";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"ff5c01e1";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"004301e1";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"27000524";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"82006b18";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"4afe2a08";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"17003304";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"ff7e01e1";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"015f01e1";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"5c01bf08";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"ef000904";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"ff5d01e1";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"ff9c01e1";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"0b006504";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"00d401e1";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"ffa701e1";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"2cff8808";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"feff8b04";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"ffa301e1";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"01ea01e1";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"ff7401e1";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"9eff4520";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"edff5010";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"3d002408";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"c3ff6604";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"00da01e1";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"ff6901e1";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"6bfeb804";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"ffa001e1";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"024801e1";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"aefe1d08";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"8b000204";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"01fc01e1";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"ff9801e1";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"beff4d04";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"009201e1";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"ff7d01e1";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"38fe9708";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"68ff2204";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"ff7401e1";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"018301e1";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"55010708";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"3d009a04";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"ff6401e1";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"000601e1";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"005f01e1";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"f5ff873c";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"15001020";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"c800260c";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"8c008f04";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"ff5c0305";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"b3ff4304";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"ff7d0305";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"011c0305";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"29ff3b0c";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"beff6c08";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"4effb004";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"019b0305";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"00280305";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"ff8b0305";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"59fe7504";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"00450305";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"ff6b0305";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"d000950c";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"1effc904";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"ff6a0305";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"62ff0804";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"016c0305";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"ffaa0305";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"27000c08";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"2a004604";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"ff8a0305";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"00cb0305";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"7affb904";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"01e20305";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"00200305";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"4afeda38";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"b7ff341c";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"2cff9210";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"a0fecb08";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"b6ff5a04";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"ffd40305";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"017c0305";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"b1feac04";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"00450305";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"ff750305";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"7efe1008";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"a9ff9a04";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"ff990305";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"01530305";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"ff620305";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"98ff8510";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"3d00b108";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"7f006404";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"ff680305";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"00710305";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"05008104";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"ff920305";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"016c0305";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"36fff308";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"9a000104";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"ff660305";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"006b0305";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"01e30305";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"14fdd108";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"71ff5204";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"ff7e0305";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"01200305";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"27010e10";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"7200d108";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"d0019704";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"ff640305";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"fff30305";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"29004f04";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"ff710305";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"015b0305";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"9dff6804";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"01520305";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"ff790305";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"f5ff8734";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"77fee924";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"e6ffe418";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"73ffec0c";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"43feec04";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"00dd0431";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"c3ffb404";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"002b0431";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"ff700431";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"f1ff6804";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"ff950431";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"5c00bb04";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"016e0431";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"ffa10431";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"c1ff4604";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"ff6a0431";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"09ff5504";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"00f10431";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"ffa40431";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"1900060c";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"e7000804";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"ff5f0431";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"40ffcf04";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"00c30431";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"ff950431";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"00ba0431";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"4afeda38";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"b7ff341c";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"2cff9210";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"afff6708";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"59ff8a04";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"ffe30431";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"01a20431";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"66002604";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"ff6d0431";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"00b20431";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"7efe1008";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"7cffb104";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"ff9e0431";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"011a0431";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"ff660431";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"98ff8510";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"3d00b108";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"7f006404";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"ff6d0431";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"00650431";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"34fffa04";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"01410431";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"ff980431";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"36fff308";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"9a000104";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"ff6a0431";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"00600431";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"016e0431";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"2500a018";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"1cfe6808";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"f1ffce04";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"ff970431";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"00db0431";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"23fe8e08";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"0800bf04";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"ff950431";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"00d20431";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"e7003d04";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"ff630431";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"ffbc0431";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"02fe0004";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"00c70431";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"92fe9a08";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"e4feea04";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"ffa60431";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"01bc0431";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"0600fd04";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"ff6a0431";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"00a40431";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"f5ff8738";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"1500101c";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"c800260c";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"8c008f04";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"ff620545";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"e5ff0b04";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"ff890545";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"00d40545";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"c800500c";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"e6ffd308";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"14fed204";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"fff00545";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"010a0545";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"ff940545";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"ff770545";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"a7ffb818";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"f1ff6908";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"6afff904";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"ff900545";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"00250545";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"0b000d08";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"25008d04";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"ff9b0545";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"00ab0545";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"44004c04";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"01540545";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"00390545";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"ff7f0545";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"27000520";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"82006b14";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"4afe2a08";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"52fefe04";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"00e60545";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"ff950545";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"5c01bf08";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"ef000904";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"ff690545";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"ffc50545";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"00730545";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"2cff8808";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"84ffd004";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"00150545";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"013c0545";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"ff870545";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"68ff1d18";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"adfec608";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"4afed204";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"01680545";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"ff9b0545";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"5aff9308";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"a1ffa304";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"ffa10545";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"01860545";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"65007e04";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"ff730545";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"00600545";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"eaff7110";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"feff9608";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"b3feb604";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"00d40545";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"ff6d0545";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"1dff2204";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"01530545";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"ffbc0545";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"98fe3704";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"00ce0545";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"4efe7504";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"00360545";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"ff620545";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"f5ff8738";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"77fee928";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"e5fefd14";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"8dfdd408";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"deffc104";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"00f50679";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"00130679";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"61fed108";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"3eff5e04";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"00a70679";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"ffa80679";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"ff6a0679";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"85ff4f04";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"ff9f0679";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"50ff4708";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"9cff5c04";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"007a0679";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"ffa30679";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"e6fffd04";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"01320679";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"00000679";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"1900060c";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"e7000804";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"ff650679";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"c5ff0804";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"00980679";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"ffa00679";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"00990679";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"4afeda30";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"b7ff761c";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"3bff8810";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"d600c608";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"35ffba04";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"ff870679";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"00650679";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"1dff7504";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"01350679";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"ff900679";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"4dfe5304";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"ff7a0679";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"8c002304";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"01520679";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"ff8b0679";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"8100480c";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"25ff3104";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"00800679";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"aefe2504";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"00170679";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"ff680679";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"3fffe104";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"015d0679";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"ff9c0679";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"2500a018";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"1cfe6808";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"a4ffac04";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"ffa20679";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"00da0679";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"ac00ee08";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"29005604";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"ff680679";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"ffca0679";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"35fef904";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"ffa00679";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"00d60679";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"14feb610";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"d1ff3508";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"3a000c04";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"ff6c0679";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"00af0679";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"cbffc804";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"ffc30679";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"01ae0679";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"3b001008";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"b1fe6b04";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"00390679";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"ff630679";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"00ae0679";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"27000534";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"82006b28";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"effff310";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"5c01bf0c";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"4afe1204";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"004f0795";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"c4006904";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"ff710795";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"000c0795";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"00780795";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"9a006b10";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"3d005808";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"4afe7f04";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"00210795";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"ff680795";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"9cff4e04";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"00eb0795";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"ffa70795";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"9a007b04";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"01c00795";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"ffa90795";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"a2ffa908";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"79ff2a04";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"001e0795";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"01020795";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"ff920795";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"15ffa124";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"94febe08";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"c3ffb304";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"011c0795";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"ff9d0795";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"b3fe840c";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"96ff1308";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"6e003004";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"01420795";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"000a0795";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"ff8a0795";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"b2005c08";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"32ffc204";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"ff630795";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"fffd0795";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"71ff8304";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"ff830795";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"01400795";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"1dff221c";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"beff4d0c";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"6e004c04";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"fffe0795";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"efff8804";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"01860795";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"00680795";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"d1ff5108";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"2cff1a04";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"009e0795";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"ffa50795";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"75fff504";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"ff890795";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"00ef0795";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"3d005210";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"c9004708";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"3fff9404";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"fff10795";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"ff650795";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"66ffe304";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"00e90795";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"ff8d0795";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"4aff0508";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"4dfe9f04";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"000c0795";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"01370795";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"ff9e0795";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"27000544";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"29ff7934";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"c1fee318";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"c300ac10";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"1f008008";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"90fe7104";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"008208e9";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"ff6708e9";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"29ff5504";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"ff7608e9";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"00d108e9";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"27ffd704";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"ffa908e9";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"00fe08e9";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"85ff940c";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"fbff1308";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"acfff004";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"00ce08e9";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"ffa808e9";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"ff6908e9";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"59001508";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"62ff3004";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"007408e9";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"ff6f08e9";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"cbffca04";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"ffe508e9";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"01c408e9";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"7200d108";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"c5febc04";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"001f08e9";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"ff6108e9";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"55ffc904";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"ffa708e9";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"00de08e9";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"15ffa128";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"79fedc10";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"f5ffac08";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"e5fea504";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"011e08e9";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"ffe708e9";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"28fe2504";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"00ab08e9";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"ff7408e9";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"2500a908";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"56fe8004";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"002d08e9";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"ff6308e9";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"48003f08";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"f2018804";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"001e08e9";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"ff8308e9";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"4bfef104";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"001608e9";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"013908e9";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"1dff2220";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"42ff8810";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"feff5208";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"b2ff4804";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"007d08e9";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"ff7808e9";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"93ff2404";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"ffbb08e9";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"00c408e9";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"70fe4608";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"1cff6c04";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"010d08e9";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"000b08e9";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"1000d904";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"ff6d08e9";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"003108e9";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"2600f210";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"3d007c08";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"2ffeaa04";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"fff308e9";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"ff6708e9";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"85003504";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"002408e9";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"00b108e9";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"aafef108";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"17ffff04";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"004108e9";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"011708e9";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"43ffa404";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"ff9208e9";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"002c08e9";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"b8ff8668";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"15ffab34";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"dbff8618";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"4fffa00c";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"4afe6a08";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"26005f04";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"00c90a0d";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"00180a0d";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"ff700a0d";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"2bfff904";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"ffaa0a0d";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"17ffcd04";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"01b60a0d";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"00250a0d";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"78ff3710";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"c1feed08";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"5affb904";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"00cf0a0d";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"ff690a0d";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"46ff5204";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"ff850a0d";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"00e90a0d";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"e5ff8108";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"adfee004";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"ffe80a0d";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"ff630a0d";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"00360a0d";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"98ff321c";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"41ffab10";
		wait for Clk_period;
		Addr <=  "0001001010111";
		Trees_din <= x"d000df08";
		wait for Clk_period;
		Addr <=  "0001001011000";
		Trees_din <= x"a3fef104";
		wait for Clk_period;
		Addr <=  "0001001011001";
		Trees_din <= x"00150a0d";
		wait for Clk_period;
		Addr <=  "0001001011010";
		Trees_din <= x"ff700a0d";
		wait for Clk_period;
		Addr <=  "0001001011011";
		Trees_din <= x"adff0504";
		wait for Clk_period;
		Addr <=  "0001001011100";
		Trees_din <= x"010c0a0d";
		wait for Clk_period;
		Addr <=  "0001001011101";
		Trees_din <= x"ffe90a0d";
		wait for Clk_period;
		Addr <=  "0001001011110";
		Trees_din <= x"51ffd704";
		wait for Clk_period;
		Addr <=  "0001001011111";
		Trees_din <= x"01f00a0d";
		wait for Clk_period;
		Addr <=  "0001001100000";
		Trees_din <= x"88003e04";
		wait for Clk_period;
		Addr <=  "0001001100001";
		Trees_din <= x"ffa70a0d";
		wait for Clk_period;
		Addr <=  "0001001100010";
		Trees_din <= x"008c0a0d";
		wait for Clk_period;
		Addr <=  "0001001100011";
		Trees_din <= x"a2ffc010";
		wait for Clk_period;
		Addr <=  "0001001100100";
		Trees_din <= x"29ffbc08";
		wait for Clk_period;
		Addr <=  "0001001100101";
		Trees_din <= x"2dff1604";
		wait for Clk_period;
		Addr <=  "0001001100110";
		Trees_din <= x"00ef0a0d";
		wait for Clk_period;
		Addr <=  "0001001100111";
		Trees_din <= x"00170a0d";
		wait for Clk_period;
		Addr <=  "0001001101000";
		Trees_din <= x"7eff0004";
		wait for Clk_period;
		Addr <=  "0001001101001";
		Trees_din <= x"ff8e0a0d";
		wait for Clk_period;
		Addr <=  "0001001101010";
		Trees_din <= x"00320a0d";
		wait for Clk_period;
		Addr <=  "0001001101011";
		Trees_din <= x"11ffd104";
		wait for Clk_period;
		Addr <=  "0001001101100";
		Trees_din <= x"ff760a0d";
		wait for Clk_period;
		Addr <=  "0001001101101";
		Trees_din <= x"00480a0d";
		wait for Clk_period;
		Addr <=  "0001001101110";
		Trees_din <= x"1c001e20";
		wait for Clk_period;
		Addr <=  "0001001101111";
		Trees_din <= x"bdfee608";
		wait for Clk_period;
		Addr <=  "0001001110000";
		Trees_din <= x"9bff0004";
		wait for Clk_period;
		Addr <=  "0001001110001";
		Trees_din <= x"01260a0d";
		wait for Clk_period;
		Addr <=  "0001001110010";
		Trees_din <= x"ff910a0d";
		wait for Clk_period;
		Addr <=  "0001001110011";
		Trees_din <= x"82006b10";
		wait for Clk_period;
		Addr <=  "0001001110100";
		Trees_din <= x"0b010208";
		wait for Clk_period;
		Addr <=  "0001001110101";
		Trees_din <= x"b4004a04";
		wait for Clk_period;
		Addr <=  "0001001110110";
		Trees_din <= x"ff6a0a0d";
		wait for Clk_period;
		Addr <=  "0001001110111";
		Trees_din <= x"002f0a0d";
		wait for Clk_period;
		Addr <=  "0001001111000";
		Trees_din <= x"f9ff6604";
		wait for Clk_period;
		Addr <=  "0001001111001";
		Trees_din <= x"ff9c0a0d";
		wait for Clk_period;
		Addr <=  "0001001111010";
		Trees_din <= x"009f0a0d";
		wait for Clk_period;
		Addr <=  "0001001111011";
		Trees_din <= x"0b003704";
		wait for Clk_period;
		Addr <=  "0001001111100";
		Trees_din <= x"ffa70a0d";
		wait for Clk_period;
		Addr <=  "0001001111101";
		Trees_din <= x"00920a0d";
		wait for Clk_period;
		Addr <=  "0001001111110";
		Trees_din <= x"77fed608";
		wait for Clk_period;
		Addr <=  "0001001111111";
		Trees_din <= x"96fee604";
		wait for Clk_period;
		Addr <=  "0001010000000";
		Trees_din <= x"00c50a0d";
		wait for Clk_period;
		Addr <=  "0001010000001";
		Trees_din <= x"00210a0d";
		wait for Clk_period;
		Addr <=  "0001010000010";
		Trees_din <= x"ff900a0d";
		wait for Clk_period;
		Addr <=  "0001010000011";
		Trees_din <= x"27000540";
		wait for Clk_period;
		Addr <=  "0001010000100";
		Trees_din <= x"29ff7930";
		wait for Clk_period;
		Addr <=  "0001010000101";
		Trees_din <= x"25001910";
		wait for Clk_period;
		Addr <=  "0001010000110";
		Trees_din <= x"78fef208";
		wait for Clk_period;
		Addr <=  "0001010000111";
		Trees_din <= x"2dff2104";
		wait for Clk_period;
		Addr <=  "0001010001000";
		Trees_din <= x"ff8f0b29";
		wait for Clk_period;
		Addr <=  "0001010001001";
		Trees_din <= x"01410b29";
		wait for Clk_period;
		Addr <=  "0001010001010";
		Trees_din <= x"ee00e904";
		wait for Clk_period;
		Addr <=  "0001010001011";
		Trees_din <= x"ff650b29";
		wait for Clk_period;
		Addr <=  "0001010001100";
		Trees_din <= x"003a0b29";
		wait for Clk_period;
		Addr <=  "0001010001101";
		Trees_din <= x"66ffe510";
		wait for Clk_period;
		Addr <=  "0001010001110";
		Trees_din <= x"da004908";
		wait for Clk_period;
		Addr <=  "0001010001111";
		Trees_din <= x"82008e04";
		wait for Clk_period;
		Addr <=  "0001010010000";
		Trees_din <= x"ff680b29";
		wait for Clk_period;
		Addr <=  "0001010010001";
		Trees_din <= x"00720b29";
		wait for Clk_period;
		Addr <=  "0001010010010";
		Trees_din <= x"c1fee704";
		wait for Clk_period;
		Addr <=  "0001010010011";
		Trees_din <= x"ffa10b29";
		wait for Clk_period;
		Addr <=  "0001010010100";
		Trees_din <= x"00e20b29";
		wait for Clk_period;
		Addr <=  "0001010010101";
		Trees_din <= x"3cff0008";
		wait for Clk_period;
		Addr <=  "0001010010110";
		Trees_din <= x"32fee204";
		wait for Clk_period;
		Addr <=  "0001010010111";
		Trees_din <= x"00d30b29";
		wait for Clk_period;
		Addr <=  "0001010011000";
		Trees_din <= x"ffb80b29";
		wait for Clk_period;
		Addr <=  "0001010011001";
		Trees_din <= x"adfeed04";
		wait for Clk_period;
		Addr <=  "0001010011010";
		Trees_din <= x"00da0b29";
		wait for Clk_period;
		Addr <=  "0001010011011";
		Trees_din <= x"ff960b29";
		wait for Clk_period;
		Addr <=  "0001010011100";
		Trees_din <= x"7200d108";
		wait for Clk_period;
		Addr <=  "0001010011101";
		Trees_din <= x"84fe9e04";
		wait for Clk_period;
		Addr <=  "0001010011110";
		Trees_din <= x"000f0b29";
		wait for Clk_period;
		Addr <=  "0001010011111";
		Trees_din <= x"ff640b29";
		wait for Clk_period;
		Addr <=  "0001010100000";
		Trees_din <= x"5eff8304";
		wait for Clk_period;
		Addr <=  "0001010100001";
		Trees_din <= x"00d80b29";
		wait for Clk_period;
		Addr <=  "0001010100010";
		Trees_din <= x"ffa80b29";
		wait for Clk_period;
		Addr <=  "0001010100011";
		Trees_din <= x"beff4d14";
		wait for Clk_period;
		Addr <=  "0001010100100";
		Trees_din <= x"baff7304";
		wait for Clk_period;
		Addr <=  "0001010100101";
		Trees_din <= x"ff9f0b29";
		wait for Clk_period;
		Addr <=  "0001010100110";
		Trees_din <= x"15ffbe08";
		wait for Clk_period;
		Addr <=  "0001010100111";
		Trees_din <= x"89ff6504";
		wait for Clk_period;
		Addr <=  "0001010101000";
		Trees_din <= x"00ab0b29";
		wait for Clk_period;
		Addr <=  "0001010101001";
		Trees_din <= x"ff990b29";
		wait for Clk_period;
		Addr <=  "0001010101010";
		Trees_din <= x"eaff9a04";
		wait for Clk_period;
		Addr <=  "0001010101011";
		Trees_din <= x"01050b29";
		wait for Clk_period;
		Addr <=  "0001010101100";
		Trees_din <= x"00340b29";
		wait for Clk_period;
		Addr <=  "0001010101101";
		Trees_din <= x"9eff3b1c";
		wait for Clk_period;
		Addr <=  "0001010101110";
		Trees_din <= x"fafee70c";
		wait for Clk_period;
		Addr <=  "0001010101111";
		Trees_din <= x"e7ffea08";
		wait for Clk_period;
		Addr <=  "0001010110000";
		Trees_din <= x"45ff1b04";
		wait for Clk_period;
		Addr <=  "0001010110001";
		Trees_din <= x"ff9c0b29";
		wait for Clk_period;
		Addr <=  "0001010110010";
		Trees_din <= x"00a00b29";
		wait for Clk_period;
		Addr <=  "0001010110011";
		Trees_din <= x"01fa0b29";
		wait for Clk_period;
		Addr <=  "0001010110100";
		Trees_din <= x"b7ff8a08";
		wait for Clk_period;
		Addr <=  "0001010110101";
		Trees_din <= x"46feed04";
		wait for Clk_period;
		Addr <=  "0001010110110";
		Trees_din <= x"ffa70b29";
		wait for Clk_period;
		Addr <=  "0001010110111";
		Trees_din <= x"00790b29";
		wait for Clk_period;
		Addr <=  "0001010111000";
		Trees_din <= x"85fee604";
		wait for Clk_period;
		Addr <=  "0001010111001";
		Trees_din <= x"00930b29";
		wait for Clk_period;
		Addr <=  "0001010111010";
		Trees_din <= x"ff6c0b29";
		wait for Clk_period;
		Addr <=  "0001010111011";
		Trees_din <= x"1eff0210";
		wait for Clk_period;
		Addr <=  "0001010111100";
		Trees_din <= x"2b005b08";
		wait for Clk_period;
		Addr <=  "0001010111101";
		Trees_din <= x"ecffac04";
		wait for Clk_period;
		Addr <=  "0001010111110";
		Trees_din <= x"00750b29";
		wait for Clk_period;
		Addr <=  "0001010111111";
		Trees_din <= x"ff930b29";
		wait for Clk_period;
		Addr <=  "0001011000000";
		Trees_din <= x"1cff0504";
		wait for Clk_period;
		Addr <=  "0001011000001";
		Trees_din <= x"010b0b29";
		wait for Clk_period;
		Addr <=  "0001011000010";
		Trees_din <= x"00260b29";
		wait for Clk_period;
		Addr <=  "0001011000011";
		Trees_din <= x"bbffbb08";
		wait for Clk_period;
		Addr <=  "0001011000100";
		Trees_din <= x"54010704";
		wait for Clk_period;
		Addr <=  "0001011000101";
		Trees_din <= x"ff6e0b29";
		wait for Clk_period;
		Addr <=  "0001011000110";
		Trees_din <= x"00020b29";
		wait for Clk_period;
		Addr <=  "0001011000111";
		Trees_din <= x"a3ff3704";
		wait for Clk_period;
		Addr <=  "0001011001000";
		Trees_din <= x"00770b29";
		wait for Clk_period;
		Addr <=  "0001011001001";
		Trees_din <= x"ff950b29";
		wait for Clk_period;
		Addr <=  "0001011001010";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0001011001011";
		Trees_din <= x"42ff895c";
		wait for Clk_period;
		Addr <=  "0001011001100";
		Trees_din <= x"0bffdb28";
		wait for Clk_period;
		Addr <=  "0001011001101";
		Trees_din <= x"23ff1114";
		wait for Clk_period;
		Addr <=  "0001011001110";
		Trees_din <= x"15ffac08";
		wait for Clk_period;
		Addr <=  "0001011001111";
		Trees_din <= x"c6feaa04";
		wait for Clk_period;
		Addr <=  "0001011010000";
		Trees_din <= x"00790c49";
		wait for Clk_period;
		Addr <=  "0001011010001";
		Trees_din <= x"ff780c49";
		wait for Clk_period;
		Addr <=  "0001011010010";
		Trees_din <= x"b5fee208";
		wait for Clk_period;
		Addr <=  "0001011010011";
		Trees_din <= x"5dffcc04";
		wait for Clk_period;
		Addr <=  "0001011010100";
		Trees_din <= x"014b0c49";
		wait for Clk_period;
		Addr <=  "0001011010101";
		Trees_din <= x"fff40c49";
		wait for Clk_period;
		Addr <=  "0001011010110";
		Trees_din <= x"ffa20c49";
		wait for Clk_period;
		Addr <=  "0001011010111";
		Trees_din <= x"7500f00c";
		wait for Clk_period;
		Addr <=  "0001011011000";
		Trees_din <= x"d0019708";
		wait for Clk_period;
		Addr <=  "0001011011001";
		Trees_din <= x"02fe0504";
		wait for Clk_period;
		Addr <=  "0001011011010";
		Trees_din <= x"00450c49";
		wait for Clk_period;
		Addr <=  "0001011011011";
		Trees_din <= x"ff700c49";
		wait for Clk_period;
		Addr <=  "0001011011100";
		Trees_din <= x"00a80c49";
		wait for Clk_period;
		Addr <=  "0001011011101";
		Trees_din <= x"72005504";
		wait for Clk_period;
		Addr <=  "0001011011110";
		Trees_din <= x"ffa70c49";
		wait for Clk_period;
		Addr <=  "0001011011111";
		Trees_din <= x"01180c49";
		wait for Clk_period;
		Addr <=  "0001011100000";
		Trees_din <= x"46fef118";
		wait for Clk_period;
		Addr <=  "0001011100001";
		Trees_din <= x"2ffefe0c";
		wait for Clk_period;
		Addr <=  "0001011100010";
		Trees_din <= x"9eff5c08";
		wait for Clk_period;
		Addr <=  "0001011100011";
		Trees_din <= x"d9ffd204";
		wait for Clk_period;
		Addr <=  "0001011100100";
		Trees_din <= x"ffe80c49";
		wait for Clk_period;
		Addr <=  "0001011100101";
		Trees_din <= x"011b0c49";
		wait for Clk_period;
		Addr <=  "0001011100110";
		Trees_din <= x"ff960c49";
		wait for Clk_period;
		Addr <=  "0001011100111";
		Trees_din <= x"33fe1204";
		wait for Clk_period;
		Addr <=  "0001011101000";
		Trees_din <= x"00730c49";
		wait for Clk_period;
		Addr <=  "0001011101001";
		Trees_din <= x"7f006404";
		wait for Clk_period;
		Addr <=  "0001011101010";
		Trees_din <= x"ff6f0c49";
		wait for Clk_period;
		Addr <=  "0001011101011";
		Trees_din <= x"004a0c49";
		wait for Clk_period;
		Addr <=  "0001011101100";
		Trees_din <= x"a2ffc910";
		wait for Clk_period;
		Addr <=  "0001011101101";
		Trees_din <= x"d4ff2b08";
		wait for Clk_period;
		Addr <=  "0001011101110";
		Trees_din <= x"99fea504";
		wait for Clk_period;
		Addr <=  "0001011101111";
		Trees_din <= x"00470c49";
		wait for Clk_period;
		Addr <=  "0001011110000";
		Trees_din <= x"ff7d0c49";
		wait for Clk_period;
		Addr <=  "0001011110001";
		Trees_din <= x"13007604";
		wait for Clk_period;
		Addr <=  "0001011110010";
		Trees_din <= x"ff930c49";
		wait for Clk_period;
		Addr <=  "0001011110011";
		Trees_din <= x"00c10c49";
		wait for Clk_period;
		Addr <=  "0001011110100";
		Trees_din <= x"54008904";
		wait for Clk_period;
		Addr <=  "0001011110101";
		Trees_din <= x"ff730c49";
		wait for Clk_period;
		Addr <=  "0001011110110";
		Trees_din <= x"e7ff5304";
		wait for Clk_period;
		Addr <=  "0001011110111";
		Trees_din <= x"00cc0c49";
		wait for Clk_period;
		Addr <=  "0001011111000";
		Trees_din <= x"ff9a0c49";
		wait for Clk_period;
		Addr <=  "0001011111001";
		Trees_din <= x"4afe780c";
		wait for Clk_period;
		Addr <=  "0001011111010";
		Trees_din <= x"e6ff8b08";
		wait for Clk_period;
		Addr <=  "0001011111011";
		Trees_din <= x"dcffea04";
		wait for Clk_period;
		Addr <=  "0001011111100";
		Trees_din <= x"ffe50c49";
		wait for Clk_period;
		Addr <=  "0001011111101";
		Trees_din <= x"01370c49";
		wait for Clk_period;
		Addr <=  "0001011111110";
		Trees_din <= x"ff8a0c49";
		wait for Clk_period;
		Addr <=  "0001011111111";
		Trees_din <= x"adff3318";
		wait for Clk_period;
		Addr <=  "0001100000000";
		Trees_din <= x"c7fea010";
		wait for Clk_period;
		Addr <=  "0001100000001";
		Trees_din <= x"9eff3d08";
		wait for Clk_period;
		Addr <=  "0001100000010";
		Trees_din <= x"dfff5a04";
		wait for Clk_period;
		Addr <=  "0001100000011";
		Trees_din <= x"00f20c49";
		wait for Clk_period;
		Addr <=  "0001100000100";
		Trees_din <= x"ffef0c49";
		wait for Clk_period;
		Addr <=  "0001100000101";
		Trees_din <= x"7bfe7f04";
		wait for Clk_period;
		Addr <=  "0001100000110";
		Trees_din <= x"001e0c49";
		wait for Clk_period;
		Addr <=  "0001100000111";
		Trees_din <= x"ff8d0c49";
		wait for Clk_period;
		Addr <=  "0001100001000";
		Trees_din <= x"5ffe6804";
		wait for Clk_period;
		Addr <=  "0001100001001";
		Trees_din <= x"00200c49";
		wait for Clk_period;
		Addr <=  "0001100001010";
		Trees_din <= x"ff700c49";
		wait for Clk_period;
		Addr <=  "0001100001011";
		Trees_din <= x"73006f08";
		wait for Clk_period;
		Addr <=  "0001100001100";
		Trees_din <= x"25011c04";
		wait for Clk_period;
		Addr <=  "0001100001101";
		Trees_din <= x"ff640c49";
		wait for Clk_period;
		Addr <=  "0001100001110";
		Trees_din <= x"00130c49";
		wait for Clk_period;
		Addr <=  "0001100001111";
		Trees_din <= x"fdffef04";
		wait for Clk_period;
		Addr <=  "0001100010000";
		Trees_din <= x"ff820c49";
		wait for Clk_period;
		Addr <=  "0001100010001";
		Trees_din <= x"00c10c49";
		wait for Clk_period;
		Addr <=  "0001100010010";
		Trees_din <= x"b8ff866c";
		wait for Clk_period;
		Addr <=  "0001100010011";
		Trees_din <= x"15ffab34";
		wait for Clk_period;
		Addr <=  "0001100010100";
		Trees_din <= x"dbff8618";
		wait for Clk_period;
		Addr <=  "0001100010101";
		Trees_din <= x"4fffa00c";
		wait for Clk_period;
		Addr <=  "0001100010110";
		Trees_din <= x"4afe6a08";
		wait for Clk_period;
		Addr <=  "0001100010111";
		Trees_din <= x"55ff8d04";
		wait for Clk_period;
		Addr <=  "0001100011000";
		Trees_din <= x"00ae0d6d";
		wait for Clk_period;
		Addr <=  "0001100011001";
		Trees_din <= x"000a0d6d";
		wait for Clk_period;
		Addr <=  "0001100011010";
		Trees_din <= x"ff7a0d6d";
		wait for Clk_period;
		Addr <=  "0001100011011";
		Trees_din <= x"68fef204";
		wait for Clk_period;
		Addr <=  "0001100011100";
		Trees_din <= x"ffde0d6d";
		wait for Clk_period;
		Addr <=  "0001100011101";
		Trees_din <= x"29ff2704";
		wait for Clk_period;
		Addr <=  "0001100011110";
		Trees_din <= x"01300d6d";
		wait for Clk_period;
		Addr <=  "0001100011111";
		Trees_din <= x"00610d6d";
		wait for Clk_period;
		Addr <=  "0001100100000";
		Trees_din <= x"78ff3710";
		wait for Clk_period;
		Addr <=  "0001100100001";
		Trees_din <= x"c1feed08";
		wait for Clk_period;
		Addr <=  "0001100100010";
		Trees_din <= x"5affb904";
		wait for Clk_period;
		Addr <=  "0001100100011";
		Trees_din <= x"00a40d6d";
		wait for Clk_period;
		Addr <=  "0001100100100";
		Trees_din <= x"ff6f0d6d";
		wait for Clk_period;
		Addr <=  "0001100100101";
		Trees_din <= x"46ff5204";
		wait for Clk_period;
		Addr <=  "0001100100110";
		Trees_din <= x"ff940d6d";
		wait for Clk_period;
		Addr <=  "0001100100111";
		Trees_din <= x"00b40d6d";
		wait for Clk_period;
		Addr <=  "0001100101000";
		Trees_din <= x"57fe2804";
		wait for Clk_period;
		Addr <=  "0001100101001";
		Trees_din <= x"003d0d6d";
		wait for Clk_period;
		Addr <=  "0001100101010";
		Trees_din <= x"adfee004";
		wait for Clk_period;
		Addr <=  "0001100101011";
		Trees_din <= x"ffec0d6d";
		wait for Clk_period;
		Addr <=  "0001100101100";
		Trees_din <= x"ff690d6d";
		wait for Clk_period;
		Addr <=  "0001100101101";
		Trees_din <= x"d1ff451c";
		wait for Clk_period;
		Addr <=  "0001100101110";
		Trees_din <= x"9dff1e0c";
		wait for Clk_period;
		Addr <=  "0001100101111";
		Trees_din <= x"58fed004";
		wait for Clk_period;
		Addr <=  "0001100110000";
		Trees_din <= x"ff8d0d6d";
		wait for Clk_period;
		Addr <=  "0001100110001";
		Trees_din <= x"31ff9804";
		wait for Clk_period;
		Addr <=  "0001100110010";
		Trees_din <= x"ffb10d6d";
		wait for Clk_period;
		Addr <=  "0001100110011";
		Trees_din <= x"00f60d6d";
		wait for Clk_period;
		Addr <=  "0001100110100";
		Trees_din <= x"38fe9708";
		wait for Clk_period;
		Addr <=  "0001100110101";
		Trees_din <= x"f8008d04";
		wait for Clk_period;
		Addr <=  "0001100110110";
		Trees_din <= x"fff70d6d";
		wait for Clk_period;
		Addr <=  "0001100110111";
		Trees_din <= x"00bb0d6d";
		wait for Clk_period;
		Addr <=  "0001100111000";
		Trees_din <= x"a2ff5404";
		wait for Clk_period;
		Addr <=  "0001100111001";
		Trees_din <= x"00360d6d";
		wait for Clk_period;
		Addr <=  "0001100111010";
		Trees_din <= x"ff810d6d";
		wait for Clk_period;
		Addr <=  "0001100111011";
		Trees_din <= x"99ff000c";
		wait for Clk_period;
		Addr <=  "0001100111100";
		Trees_din <= x"5fff7a08";
		wait for Clk_period;
		Addr <=  "0001100111101";
		Trees_din <= x"b1fee904";
		wait for Clk_period;
		Addr <=  "0001100111110";
		Trees_din <= x"010d0d6d";
		wait for Clk_period;
		Addr <=  "0001100111111";
		Trees_din <= x"00540d6d";
		wait for Clk_period;
		Addr <=  "0001101000000";
		Trees_din <= x"ff970d6d";
		wait for Clk_period;
		Addr <=  "0001101000001";
		Trees_din <= x"cdff8008";
		wait for Clk_period;
		Addr <=  "0001101000010";
		Trees_din <= x"7bff7304";
		wait for Clk_period;
		Addr <=  "0001101000011";
		Trees_din <= x"ffa30d6d";
		wait for Clk_period;
		Addr <=  "0001101000100";
		Trees_din <= x"00970d6d";
		wait for Clk_period;
		Addr <=  "0001101000101";
		Trees_din <= x"e7ffed04";
		wait for Clk_period;
		Addr <=  "0001101000110";
		Trees_din <= x"ff790d6d";
		wait for Clk_period;
		Addr <=  "0001101000111";
		Trees_din <= x"ffe00d6d";
		wait for Clk_period;
		Addr <=  "0001101001000";
		Trees_din <= x"bdfee608";
		wait for Clk_period;
		Addr <=  "0001101001001";
		Trees_din <= x"9bff0004";
		wait for Clk_period;
		Addr <=  "0001101001010";
		Trees_din <= x"00de0d6d";
		wait for Clk_period;
		Addr <=  "0001101001011";
		Trees_din <= x"ffa10d6d";
		wait for Clk_period;
		Addr <=  "0001101001100";
		Trees_din <= x"1c001e14";
		wait for Clk_period;
		Addr <=  "0001101001101";
		Trees_din <= x"82006b10";
		wait for Clk_period;
		Addr <=  "0001101001110";
		Trees_din <= x"0b010208";
		wait for Clk_period;
		Addr <=  "0001101001111";
		Trees_din <= x"95ffd504";
		wait for Clk_period;
		Addr <=  "0001101010000";
		Trees_din <= x"ff690d6d";
		wait for Clk_period;
		Addr <=  "0001101010001";
		Trees_din <= x"ffd30d6d";
		wait for Clk_period;
		Addr <=  "0001101010010";
		Trees_din <= x"81ffd104";
		wait for Clk_period;
		Addr <=  "0001101010011";
		Trees_din <= x"ffab0d6d";
		wait for Clk_period;
		Addr <=  "0001101010100";
		Trees_din <= x"00860d6d";
		wait for Clk_period;
		Addr <=  "0001101010101";
		Trees_din <= x"00270d6d";
		wait for Clk_period;
		Addr <=  "0001101010110";
		Trees_din <= x"77fed608";
		wait for Clk_period;
		Addr <=  "0001101010111";
		Trees_din <= x"cdff4004";
		wait for Clk_period;
		Addr <=  "0001101011000";
		Trees_din <= x"00960d6d";
		wait for Clk_period;
		Addr <=  "0001101011001";
		Trees_din <= x"001b0d6d";
		wait for Clk_period;
		Addr <=  "0001101011010";
		Trees_din <= x"ffa20d6d";
		wait for Clk_period;
		Addr <=  "0001101011011";
		Trees_din <= x"42ffa550";
		wait for Clk_period;
		Addr <=  "0001101011100";
		Trees_din <= x"58fea918";
		wait for Clk_period;
		Addr <=  "0001101011101";
		Trees_din <= x"3000460c";
		wait for Clk_period;
		Addr <=  "0001101011110";
		Trees_din <= x"d0016908";
		wait for Clk_period;
		Addr <=  "0001101011111";
		Trees_din <= x"f3ffb604";
		wait for Clk_period;
		Addr <=  "0001101100000";
		Trees_din <= x"ff680e59";
		wait for Clk_period;
		Addr <=  "0001101100001";
		Trees_din <= x"001d0e59";
		wait for Clk_period;
		Addr <=  "0001101100010";
		Trees_din <= x"00400e59";
		wait for Clk_period;
		Addr <=  "0001101100011";
		Trees_din <= x"e6000c08";
		wait for Clk_period;
		Addr <=  "0001101100100";
		Trees_din <= x"7fffc904";
		wait for Clk_period;
		Addr <=  "0001101100101";
		Trees_din <= x"ff940e59";
		wait for Clk_period;
		Addr <=  "0001101100110";
		Trees_din <= x"fff60e59";
		wait for Clk_period;
		Addr <=  "0001101100111";
		Trees_din <= x"00c00e59";
		wait for Clk_period;
		Addr <=  "0001101101000";
		Trees_din <= x"9eff4518";
		wait for Clk_period;
		Addr <=  "0001101101001";
		Trees_din <= x"b4ff4410";
		wait for Clk_period;
		Addr <=  "0001101101010";
		Trees_din <= x"e7000808";
		wait for Clk_period;
		Addr <=  "0001101101011";
		Trees_din <= x"78ffa904";
		wait for Clk_period;
		Addr <=  "0001101101100";
		Trees_din <= x"00630e59";
		wait for Clk_period;
		Addr <=  "0001101101101";
		Trees_din <= x"ffaa0e59";
		wait for Clk_period;
		Addr <=  "0001101101110";
		Trees_din <= x"ecffc404";
		wait for Clk_period;
		Addr <=  "0001101101111";
		Trees_din <= x"01560e59";
		wait for Clk_period;
		Addr <=  "0001101110000";
		Trees_din <= x"00140e59";
		wait for Clk_period;
		Addr <=  "0001101110001";
		Trees_din <= x"a1fe9304";
		wait for Clk_period;
		Addr <=  "0001101110010";
		Trees_din <= x"00530e59";
		wait for Clk_period;
		Addr <=  "0001101110011";
		Trees_din <= x"ff770e59";
		wait for Clk_period;
		Addr <=  "0001101110100";
		Trees_din <= x"0bfff310";
		wait for Clk_period;
		Addr <=  "0001101110101";
		Trees_din <= x"09004908";
		wait for Clk_period;
		Addr <=  "0001101110110";
		Trees_din <= x"e0ffed04";
		wait for Clk_period;
		Addr <=  "0001101110111";
		Trees_din <= x"ff790e59";
		wait for Clk_period;
		Addr <=  "0001101111000";
		Trees_din <= x"00420e59";
		wait for Clk_period;
		Addr <=  "0001101111001";
		Trees_din <= x"c4ff3d04";
		wait for Clk_period;
		Addr <=  "0001101111010";
		Trees_din <= x"ffa60e59";
		wait for Clk_period;
		Addr <=  "0001101111011";
		Trees_din <= x"01160e59";
		wait for Clk_period;
		Addr <=  "0001101111100";
		Trees_din <= x"f8008b08";
		wait for Clk_period;
		Addr <=  "0001101111101";
		Trees_din <= x"23ff5b04";
		wait for Clk_period;
		Addr <=  "0001101111110";
		Trees_din <= x"00520e59";
		wait for Clk_period;
		Addr <=  "0001101111111";
		Trees_din <= x"ff980e59";
		wait for Clk_period;
		Addr <=  "0001110000000";
		Trees_din <= x"b1ff0e04";
		wait for Clk_period;
		Addr <=  "0001110000001";
		Trees_din <= x"00d10e59";
		wait for Clk_period;
		Addr <=  "0001110000010";
		Trees_din <= x"ffc00e59";
		wait for Clk_period;
		Addr <=  "0001110000011";
		Trees_din <= x"14fe4c10";
		wait for Clk_period;
		Addr <=  "0001110000100";
		Trees_din <= x"aefe7108";
		wait for Clk_period;
		Addr <=  "0001110000101";
		Trees_din <= x"cefff404";
		wait for Clk_period;
		Addr <=  "0001110000110";
		Trees_din <= x"00b90e59";
		wait for Clk_period;
		Addr <=  "0001110000111";
		Trees_din <= x"00000e59";
		wait for Clk_period;
		Addr <=  "0001110001000";
		Trees_din <= x"93fef404";
		wait for Clk_period;
		Addr <=  "0001110001001";
		Trees_din <= x"fff60e59";
		wait for Clk_period;
		Addr <=  "0001110001010";
		Trees_din <= x"ff940e59";
		wait for Clk_period;
		Addr <=  "0001110001011";
		Trees_din <= x"5100990c";
		wait for Clk_period;
		Addr <=  "0001110001100";
		Trees_din <= x"1700b308";
		wait for Clk_period;
		Addr <=  "0001110001101";
		Trees_din <= x"1200ef04";
		wait for Clk_period;
		Addr <=  "0001110001110";
		Trees_din <= x"ff660e59";
		wait for Clk_period;
		Addr <=  "0001110001111";
		Trees_din <= x"fffe0e59";
		wait for Clk_period;
		Addr <=  "0001110010000";
		Trees_din <= x"00010e59";
		wait for Clk_period;
		Addr <=  "0001110010001";
		Trees_din <= x"46ff2d04";
		wait for Clk_period;
		Addr <=  "0001110010010";
		Trees_din <= x"ff820e59";
		wait for Clk_period;
		Addr <=  "0001110010011";
		Trees_din <= x"46ff4304";
		wait for Clk_period;
		Addr <=  "0001110010100";
		Trees_din <= x"00a90e59";
		wait for Clk_period;
		Addr <=  "0001110010101";
		Trees_din <= x"ffad0e59";
		wait for Clk_period;
		Addr <=  "0001110010110";
		Trees_din <= x"42ffa564";
		wait for Clk_period;
		Addr <=  "0001110010111";
		Trees_din <= x"c1fed330";
		wait for Clk_period;
		Addr <=  "0001110011000";
		Trees_din <= x"7500f020";
		wait for Clk_period;
		Addr <=  "0001110011001";
		Trees_din <= x"66ffdf10";
		wait for Clk_period;
		Addr <=  "0001110011010";
		Trees_din <= x"4800b308";
		wait for Clk_period;
		Addr <=  "0001110011011";
		Trees_din <= x"f5ff6c04";
		wait for Clk_period;
		Addr <=  "0001110011100";
		Trees_din <= x"00170f65";
		wait for Clk_period;
		Addr <=  "0001110011101";
		Trees_din <= x"ff680f65";
		wait for Clk_period;
		Addr <=  "0001110011110";
		Trees_din <= x"75006504";
		wait for Clk_period;
		Addr <=  "0001110011111";
		Trees_din <= x"ffa50f65";
		wait for Clk_period;
		Addr <=  "0001110100000";
		Trees_din <= x"009f0f65";
		wait for Clk_period;
		Addr <=  "0001110100001";
		Trees_din <= x"05007208";
		wait for Clk_period;
		Addr <=  "0001110100010";
		Trees_din <= x"21003a04";
		wait for Clk_period;
		Addr <=  "0001110100011";
		Trees_din <= x"ff710f65";
		wait for Clk_period;
		Addr <=  "0001110100100";
		Trees_din <= x"00640f65";
		wait for Clk_period;
		Addr <=  "0001110100101";
		Trees_din <= x"2fff6e04";
		wait for Clk_period;
		Addr <=  "0001110100110";
		Trees_din <= x"005b0f65";
		wait for Clk_period;
		Addr <=  "0001110100111";
		Trees_din <= x"ff840f65";
		wait for Clk_period;
		Addr <=  "0001110101000";
		Trees_din <= x"9eff3d08";
		wait for Clk_period;
		Addr <=  "0001110101001";
		Trees_din <= x"01fe8704";
		wait for Clk_period;
		Addr <=  "0001110101010";
		Trees_din <= x"003f0f65";
		wait for Clk_period;
		Addr <=  "0001110101011";
		Trees_din <= x"01400f65";
		wait for Clk_period;
		Addr <=  "0001110101100";
		Trees_din <= x"45ff0204";
		wait for Clk_period;
		Addr <=  "0001110101101";
		Trees_din <= x"ffae0f65";
		wait for Clk_period;
		Addr <=  "0001110101110";
		Trees_din <= x"000f0f65";
		wait for Clk_period;
		Addr <=  "0001110101111";
		Trees_din <= x"29ff741c";
		wait for Clk_period;
		Addr <=  "0001110110000";
		Trees_din <= x"b1fee20c";
		wait for Clk_period;
		Addr <=  "0001110110001";
		Trees_din <= x"e4fe8104";
		wait for Clk_period;
		Addr <=  "0001110110010";
		Trees_din <= x"ff9b0f65";
		wait for Clk_period;
		Addr <=  "0001110110011";
		Trees_din <= x"e2ff4b04";
		wait for Clk_period;
		Addr <=  "0001110110100";
		Trees_din <= x"00680f65";
		wait for Clk_period;
		Addr <=  "0001110110101";
		Trees_din <= x"01330f65";
		wait for Clk_period;
		Addr <=  "0001110110110";
		Trees_din <= x"78ff0608";
		wait for Clk_period;
		Addr <=  "0001110110111";
		Trees_din <= x"1eff5d04";
		wait for Clk_period;
		Addr <=  "0001110111000";
		Trees_din <= x"00af0f65";
		wait for Clk_period;
		Addr <=  "0001110111001";
		Trees_din <= x"ffdb0f65";
		wait for Clk_period;
		Addr <=  "0001110111010";
		Trees_din <= x"9cfef404";
		wait for Clk_period;
		Addr <=  "0001110111011";
		Trees_din <= x"006c0f65";
		wait for Clk_period;
		Addr <=  "0001110111100";
		Trees_din <= x"ffac0f65";
		wait for Clk_period;
		Addr <=  "0001110111101";
		Trees_din <= x"29005610";
		wait for Clk_period;
		Addr <=  "0001110111110";
		Trees_din <= x"4afe7f08";
		wait for Clk_period;
		Addr <=  "0001110111111";
		Trees_din <= x"09ffe504";
		wait for Clk_period;
		Addr <=  "0001111000000";
		Trees_din <= x"00000f65";
		wait for Clk_period;
		Addr <=  "0001111000001";
		Trees_din <= x"00840f65";
		wait for Clk_period;
		Addr <=  "0001111000010";
		Trees_din <= x"95fff204";
		wait for Clk_period;
		Addr <=  "0001111000011";
		Trees_din <= x"ff6c0f65";
		wait for Clk_period;
		Addr <=  "0001111000100";
		Trees_din <= x"001d0f65";
		wait for Clk_period;
		Addr <=  "0001111000101";
		Trees_din <= x"aefecd04";
		wait for Clk_period;
		Addr <=  "0001111000110";
		Trees_din <= x"00df0f65";
		wait for Clk_period;
		Addr <=  "0001111000111";
		Trees_din <= x"ffa60f65";
		wait for Clk_period;
		Addr <=  "0001111001000";
		Trees_din <= x"4afe850c";
		wait for Clk_period;
		Addr <=  "0001111001001";
		Trees_din <= x"85ffcf04";
		wait for Clk_period;
		Addr <=  "0001111001010";
		Trees_din <= x"ff9a0f65";
		wait for Clk_period;
		Addr <=  "0001111001011";
		Trees_din <= x"82ff1204";
		wait for Clk_period;
		Addr <=  "0001111001100";
		Trees_din <= x"ffef0f65";
		wait for Clk_period;
		Addr <=  "0001111001101";
		Trees_din <= x"009c0f65";
		wait for Clk_period;
		Addr <=  "0001111001110";
		Trees_din <= x"8c00b00c";
		wait for Clk_period;
		Addr <=  "0001111001111";
		Trees_din <= x"b1fe7d08";
		wait for Clk_period;
		Addr <=  "0001111010000";
		Trees_din <= x"6c000604";
		wait for Clk_period;
		Addr <=  "0001111010001";
		Trees_din <= x"ff960f65";
		wait for Clk_period;
		Addr <=  "0001111010010";
		Trees_din <= x"006c0f65";
		wait for Clk_period;
		Addr <=  "0001111010011";
		Trees_din <= x"ff670f65";
		wait for Clk_period;
		Addr <=  "0001111010100";
		Trees_din <= x"d2fe7008";
		wait for Clk_period;
		Addr <=  "0001111010101";
		Trees_din <= x"48003304";
		wait for Clk_period;
		Addr <=  "0001111010110";
		Trees_din <= x"000f0f65";
		wait for Clk_period;
		Addr <=  "0001111010111";
		Trees_din <= x"00930f65";
		wait for Clk_period;
		Addr <=  "0001111011000";
		Trees_din <= x"ff910f65";
		wait for Clk_period;
		Addr <=  "0001111011001";
		Trees_din <= x"42ffa558";
		wait for Clk_period;
		Addr <=  "0001111011010";
		Trees_din <= x"58fea91c";
		wait for Clk_period;
		Addr <=  "0001111011011";
		Trees_din <= x"1aff1b08";
		wait for Clk_period;
		Addr <=  "0001111011100";
		Trees_din <= x"cafd9004";
		wait for Clk_period;
		Addr <=  "0001111011101";
		Trees_din <= x"00061051";
		wait for Clk_period;
		Addr <=  "0001111011110";
		Trees_din <= x"ff6b1051";
		wait for Clk_period;
		Addr <=  "0001111011111";
		Trees_din <= x"34002208";
		wait for Clk_period;
		Addr <=  "0001111100000";
		Trees_din <= x"f6fe8404";
		wait for Clk_period;
		Addr <=  "0001111100001";
		Trees_din <= x"fff01051";
		wait for Clk_period;
		Addr <=  "0001111100010";
		Trees_din <= x"ff851051";
		wait for Clk_period;
		Addr <=  "0001111100011";
		Trees_din <= x"52ff0508";
		wait for Clk_period;
		Addr <=  "0001111100100";
		Trees_din <= x"e6ffec04";
		wait for Clk_period;
		Addr <=  "0001111100101";
		Trees_din <= x"00321051";
		wait for Clk_period;
		Addr <=  "0001111100110";
		Trees_din <= x"00ff1051";
		wait for Clk_period;
		Addr <=  "0001111100111";
		Trees_din <= x"ffb11051";
		wait for Clk_period;
		Addr <=  "0001111101000";
		Trees_din <= x"b4ff1a20";
		wait for Clk_period;
		Addr <=  "0001111101001";
		Trees_din <= x"79ff1010";
		wait for Clk_period;
		Addr <=  "0001111101010";
		Trees_din <= x"46feb708";
		wait for Clk_period;
		Addr <=  "0001111101011";
		Trees_din <= x"17ff6f04";
		wait for Clk_period;
		Addr <=  "0001111101100";
		Trees_din <= x"00411051";
		wait for Clk_period;
		Addr <=  "0001111101101";
		Trees_din <= x"ff831051";
		wait for Clk_period;
		Addr <=  "0001111101110";
		Trees_din <= x"53ffea04";
		wait for Clk_period;
		Addr <=  "0001111101111";
		Trees_din <= x"00a41051";
		wait for Clk_period;
		Addr <=  "0001111110000";
		Trees_din <= x"ffa01051";
		wait for Clk_period;
		Addr <=  "0001111110001";
		Trees_din <= x"adff4208";
		wait for Clk_period;
		Addr <=  "0001111110010";
		Trees_din <= x"c3fff204";
		wait for Clk_period;
		Addr <=  "0001111110011";
		Trees_din <= x"009a1051";
		wait for Clk_period;
		Addr <=  "0001111110100";
		Trees_din <= x"ffcb1051";
		wait for Clk_period;
		Addr <=  "0001111110101";
		Trees_din <= x"c1ff0704";
		wait for Clk_period;
		Addr <=  "0001111110110";
		Trees_din <= x"ff931051";
		wait for Clk_period;
		Addr <=  "0001111110111";
		Trees_din <= x"00251051";
		wait for Clk_period;
		Addr <=  "0001111111000";
		Trees_din <= x"4400420c";
		wait for Clk_period;
		Addr <=  "0001111111001";
		Trees_din <= x"bafed604";
		wait for Clk_period;
		Addr <=  "0001111111010";
		Trees_din <= x"00701051";
		wait for Clk_period;
		Addr <=  "0001111111011";
		Trees_din <= x"b2005f04";
		wait for Clk_period;
		Addr <=  "0001111111100";
		Trees_din <= x"ff711051";
		wait for Clk_period;
		Addr <=  "0001111111101";
		Trees_din <= x"00551051";
		wait for Clk_period;
		Addr <=  "0001111111110";
		Trees_din <= x"b5fed008";
		wait for Clk_period;
		Addr <=  "0001111111111";
		Trees_din <= x"ed000504";
		wait for Clk_period;
		Addr <=  "0010000000000";
		Trees_din <= x"00051051";
		wait for Clk_period;
		Addr <=  "0010000000001";
		Trees_din <= x"00eb1051";
		wait for Clk_period;
		Addr <=  "0010000000010";
		Trees_din <= x"44008a04";
		wait for Clk_period;
		Addr <=  "0010000000011";
		Trees_din <= x"ff941051";
		wait for Clk_period;
		Addr <=  "0010000000100";
		Trees_din <= x"fff91051";
		wait for Clk_period;
		Addr <=  "0010000000101";
		Trees_din <= x"e2fea514";
		wait for Clk_period;
		Addr <=  "0010000000110";
		Trees_din <= x"aefe9f0c";
		wait for Clk_period;
		Addr <=  "0010000000111";
		Trees_din <= x"2cff3904";
		wait for Clk_period;
		Addr <=  "0010000001000";
		Trees_din <= x"00a71051";
		wait for Clk_period;
		Addr <=  "0010000001001";
		Trees_din <= x"edff5304";
		wait for Clk_period;
		Addr <=  "0010000001010";
		Trees_din <= x"003c1051";
		wait for Clk_period;
		Addr <=  "0010000001011";
		Trees_din <= x"ffb11051";
		wait for Clk_period;
		Addr <=  "0010000001100";
		Trees_din <= x"66ff9304";
		wait for Clk_period;
		Addr <=  "0010000001101";
		Trees_din <= x"ffed1051";
		wait for Clk_period;
		Addr <=  "0010000001110";
		Trees_din <= x"ff8e1051";
		wait for Clk_period;
		Addr <=  "0010000001111";
		Trees_din <= x"4afe6a04";
		wait for Clk_period;
		Addr <=  "0010000010000";
		Trees_din <= x"001a1051";
		wait for Clk_period;
		Addr <=  "0010000010001";
		Trees_din <= x"d2fe0304";
		wait for Clk_period;
		Addr <=  "0010000010010";
		Trees_din <= x"00201051";
		wait for Clk_period;
		Addr <=  "0010000010011";
		Trees_din <= x"ff681051";
		wait for Clk_period;
		Addr <=  "0010000010100";
		Trees_din <= x"b8ff8650";
		wait for Clk_period;
		Addr <=  "0010000010101";
		Trees_din <= x"15ffab28";
		wait for Clk_period;
		Addr <=  "0010000010110";
		Trees_din <= x"dbff8610";
		wait for Clk_period;
		Addr <=  "0010000010111";
		Trees_din <= x"88fff004";
		wait for Clk_period;
		Addr <=  "0010000011000";
		Trees_din <= x"ff931145";
		wait for Clk_period;
		Addr <=  "0010000011001";
		Trees_din <= x"68fec704";
		wait for Clk_period;
		Addr <=  "0010000011010";
		Trees_din <= x"ffaf1145";
		wait for Clk_period;
		Addr <=  "0010000011011";
		Trees_din <= x"f1ff7b04";
		wait for Clk_period;
		Addr <=  "0010000011100";
		Trees_din <= x"00011145";
		wait for Clk_period;
		Addr <=  "0010000011101";
		Trees_din <= x"00ac1145";
		wait for Clk_period;
		Addr <=  "0010000011110";
		Trees_din <= x"78ff370c";
		wait for Clk_period;
		Addr <=  "0010000011111";
		Trees_din <= x"46ff0304";
		wait for Clk_period;
		Addr <=  "0010000100000";
		Trees_din <= x"ff7f1145";
		wait for Clk_period;
		Addr <=  "0010000100001";
		Trees_din <= x"7dff9c04";
		wait for Clk_period;
		Addr <=  "0010000100010";
		Trees_din <= x"ff8e1145";
		wait for Clk_period;
		Addr <=  "0010000100011";
		Trees_din <= x"00761145";
		wait for Clk_period;
		Addr <=  "0010000100100";
		Trees_din <= x"e5ff8108";
		wait for Clk_period;
		Addr <=  "0010000100101";
		Trees_din <= x"adfee004";
		wait for Clk_period;
		Addr <=  "0010000100110";
		Trees_din <= x"fffa1145";
		wait for Clk_period;
		Addr <=  "0010000100111";
		Trees_din <= x"ff6a1145";
		wait for Clk_period;
		Addr <=  "0010000101000";
		Trees_din <= x"00591145";
		wait for Clk_period;
		Addr <=  "0010000101001";
		Trees_din <= x"98ff2318";
		wait for Clk_period;
		Addr <=  "0010000101010";
		Trees_din <= x"41ffab10";
		wait for Clk_period;
		Addr <=  "0010000101011";
		Trees_din <= x"04007c08";
		wait for Clk_period;
		Addr <=  "0010000101100";
		Trees_din <= x"78fe7504";
		wait for Clk_period;
		Addr <=  "0010000101101";
		Trees_din <= x"00201145";
		wait for Clk_period;
		Addr <=  "0010000101110";
		Trees_din <= x"ff791145";
		wait for Clk_period;
		Addr <=  "0010000101111";
		Trees_din <= x"fdff9304";
		wait for Clk_period;
		Addr <=  "0010000110000";
		Trees_din <= x"ffcb1145";
		wait for Clk_period;
		Addr <=  "0010000110001";
		Trees_din <= x"00661145";
		wait for Clk_period;
		Addr <=  "0010000110010";
		Trees_din <= x"51ffd704";
		wait for Clk_period;
		Addr <=  "0010000110011";
		Trees_din <= x"00ce1145";
		wait for Clk_period;
		Addr <=  "0010000110100";
		Trees_din <= x"00061145";
		wait for Clk_period;
		Addr <=  "0010000110101";
		Trees_din <= x"20005a0c";
		wait for Clk_period;
		Addr <=  "0010000110110";
		Trees_din <= x"25ffbb04";
		wait for Clk_period;
		Addr <=  "0010000110111";
		Trees_din <= x"ffa31145";
		wait for Clk_period;
		Addr <=  "0010000111000";
		Trees_din <= x"9eff7804";
		wait for Clk_period;
		Addr <=  "0010000111001";
		Trees_din <= x"00a81145";
		wait for Clk_period;
		Addr <=  "0010000111010";
		Trees_din <= x"00141145";
		wait for Clk_period;
		Addr <=  "0010000111011";
		Trees_din <= x"ffa81145";
		wait for Clk_period;
		Addr <=  "0010000111100";
		Trees_din <= x"fbff2b10";
		wait for Clk_period;
		Addr <=  "0010000111101";
		Trees_din <= x"dbffec0c";
		wait for Clk_period;
		Addr <=  "0010000111110";
		Trees_din <= x"f5fff808";
		wait for Clk_period;
		Addr <=  "0010000111111";
		Trees_din <= x"be000704";
		wait for Clk_period;
		Addr <=  "0010001000000";
		Trees_din <= x"00031145";
		wait for Clk_period;
		Addr <=  "0010001000001";
		Trees_din <= x"00d31145";
		wait for Clk_period;
		Addr <=  "0010001000010";
		Trees_din <= x"ffa91145";
		wait for Clk_period;
		Addr <=  "0010001000011";
		Trees_din <= x"ff831145";
		wait for Clk_period;
		Addr <=  "0010001000100";
		Trees_din <= x"7efe430c";
		wait for Clk_period;
		Addr <=  "0010001000101";
		Trees_din <= x"28ff8208";
		wait for Clk_period;
		Addr <=  "0010001000110";
		Trees_din <= x"03001904";
		wait for Clk_period;
		Addr <=  "0010001000111";
		Trees_din <= x"ff891145";
		wait for Clk_period;
		Addr <=  "0010001001000";
		Trees_din <= x"00191145";
		wait for Clk_period;
		Addr <=  "0010001001001";
		Trees_din <= x"00851145";
		wait for Clk_period;
		Addr <=  "0010001001010";
		Trees_din <= x"57fdfd04";
		wait for Clk_period;
		Addr <=  "0010001001011";
		Trees_din <= x"00251145";
		wait for Clk_period;
		Addr <=  "0010001001100";
		Trees_din <= x"20004304";
		wait for Clk_period;
		Addr <=  "0010001001101";
		Trees_din <= x"ff691145";
		wait for Clk_period;
		Addr <=  "0010001001110";
		Trees_din <= x"5dffeb04";
		wait for Clk_period;
		Addr <=  "0010001001111";
		Trees_din <= x"ff991145";
		wait for Clk_period;
		Addr <=  "0010001010000";
		Trees_din <= x"004b1145";
		wait for Clk_period;
		Addr <=  "0010001010001";
		Trees_din <= x"42ffa544";
		wait for Clk_period;
		Addr <=  "0010001010010";
		Trees_din <= x"58fea918";
		wait for Clk_period;
		Addr <=  "0010001010011";
		Trees_din <= x"1aff1b08";
		wait for Clk_period;
		Addr <=  "0010001010100";
		Trees_din <= x"bcffbf04";
		wait for Clk_period;
		Addr <=  "0010001010101";
		Trees_din <= x"ff6e1211";
		wait for Clk_period;
		Addr <=  "0010001010110";
		Trees_din <= x"00081211";
		wait for Clk_period;
		Addr <=  "0010001010111";
		Trees_din <= x"34002208";
		wait for Clk_period;
		Addr <=  "0010001011000";
		Trees_din <= x"f4ff3b04";
		wait for Clk_period;
		Addr <=  "0010001011001";
		Trees_din <= x"ff8e1211";
		wait for Clk_period;
		Addr <=  "0010001011010";
		Trees_din <= x"ffec1211";
		wait for Clk_period;
		Addr <=  "0010001011011";
		Trees_din <= x"e6fffb04";
		wait for Clk_period;
		Addr <=  "0010001011100";
		Trees_din <= x"fffd1211";
		wait for Clk_period;
		Addr <=  "0010001011101";
		Trees_din <= x"00c51211";
		wait for Clk_period;
		Addr <=  "0010001011110";
		Trees_din <= x"0bff850c";
		wait for Clk_period;
		Addr <=  "0010001011111";
		Trees_din <= x"ce002308";
		wait for Clk_period;
		Addr <=  "0010001100000";
		Trees_din <= x"5c00f404";
		wait for Clk_period;
		Addr <=  "0010001100001";
		Trees_din <= x"ff731211";
		wait for Clk_period;
		Addr <=  "0010001100010";
		Trees_din <= x"00091211";
		wait for Clk_period;
		Addr <=  "0010001100011";
		Trees_din <= x"00471211";
		wait for Clk_period;
		Addr <=  "0010001100100";
		Trees_din <= x"79ff1310";
		wait for Clk_period;
		Addr <=  "0010001100101";
		Trees_din <= x"d3feb608";
		wait for Clk_period;
		Addr <=  "0010001100110";
		Trees_din <= x"3d005204";
		wait for Clk_period;
		Addr <=  "0010001100111";
		Trees_din <= x"ff8e1211";
		wait for Clk_period;
		Addr <=  "0010001101000";
		Trees_din <= x"002e1211";
		wait for Clk_period;
		Addr <=  "0010001101001";
		Trees_din <= x"0fffe804";
		wait for Clk_period;
		Addr <=  "0010001101010";
		Trees_din <= x"007e1211";
		wait for Clk_period;
		Addr <=  "0010001101011";
		Trees_din <= x"ffb91211";
		wait for Clk_period;
		Addr <=  "0010001101100";
		Trees_din <= x"68fec908";
		wait for Clk_period;
		Addr <=  "0010001101101";
		Trees_din <= x"2cff6604";
		wait for Clk_period;
		Addr <=  "0010001101110";
		Trees_din <= x"00211211";
		wait for Clk_period;
		Addr <=  "0010001101111";
		Trees_din <= x"ff711211";
		wait for Clk_period;
		Addr <=  "0010001110000";
		Trees_din <= x"d1ff4504";
		wait for Clk_period;
		Addr <=  "0010001110001";
		Trees_din <= x"ffce1211";
		wait for Clk_period;
		Addr <=  "0010001110010";
		Trees_din <= x"005a1211";
		wait for Clk_period;
		Addr <=  "0010001110011";
		Trees_din <= x"14fe4c0c";
		wait for Clk_period;
		Addr <=  "0010001110100";
		Trees_din <= x"aefe7108";
		wait for Clk_period;
		Addr <=  "0010001110101";
		Trees_din <= x"d1ff5204";
		wait for Clk_period;
		Addr <=  "0010001110110";
		Trees_din <= x"00211211";
		wait for Clk_period;
		Addr <=  "0010001110111";
		Trees_din <= x"00991211";
		wait for Clk_period;
		Addr <=  "0010001111000";
		Trees_din <= x"ffbc1211";
		wait for Clk_period;
		Addr <=  "0010001111001";
		Trees_din <= x"5100990c";
		wait for Clk_period;
		Addr <=  "0010001111010";
		Trees_din <= x"7c008104";
		wait for Clk_period;
		Addr <=  "0010001111011";
		Trees_din <= x"ff6a1211";
		wait for Clk_period;
		Addr <=  "0010001111100";
		Trees_din <= x"4dfeda04";
		wait for Clk_period;
		Addr <=  "0010001111101";
		Trees_din <= x"ffa91211";
		wait for Clk_period;
		Addr <=  "0010001111110";
		Trees_din <= x"002e1211";
		wait for Clk_period;
		Addr <=  "0010001111111";
		Trees_din <= x"88000d08";
		wait for Clk_period;
		Addr <=  "0010010000000";
		Trees_din <= x"13009604";
		wait for Clk_period;
		Addr <=  "0010010000001";
		Trees_din <= x"00781211";
		wait for Clk_period;
		Addr <=  "0010010000010";
		Trees_din <= x"fff11211";
		wait for Clk_period;
		Addr <=  "0010010000011";
		Trees_din <= x"ff931211";
		wait for Clk_period;
		Addr <=  "0010010000100";
		Trees_din <= x"b8ff864c";
		wait for Clk_period;
		Addr <=  "0010010000101";
		Trees_din <= x"b4ff1a30";
		wait for Clk_period;
		Addr <=  "0010010000110";
		Trees_din <= x"78ffaf20";
		wait for Clk_period;
		Addr <=  "0010010000111";
		Trees_din <= x"9eff7810";
		wait for Clk_period;
		Addr <=  "0010010001000";
		Trees_din <= x"98feb108";
		wait for Clk_period;
		Addr <=  "0010010001001";
		Trees_din <= x"12003d04";
		wait for Clk_period;
		Addr <=  "0010010001010";
		Trees_din <= x"ff8212ed";
		wait for Clk_period;
		Addr <=  "0010010001011";
		Trees_din <= x"004712ed";
		wait for Clk_period;
		Addr <=  "0010010001100";
		Trees_din <= x"c0ff1804";
		wait for Clk_period;
		Addr <=  "0010010001101";
		Trees_din <= x"ffbb12ed";
		wait for Clk_period;
		Addr <=  "0010010001110";
		Trees_din <= x"007e12ed";
		wait for Clk_period;
		Addr <=  "0010010001111";
		Trees_din <= x"9dffe908";
		wait for Clk_period;
		Addr <=  "0010010010000";
		Trees_din <= x"91ffe804";
		wait for Clk_period;
		Addr <=  "0010010010001";
		Trees_din <= x"ff9512ed";
		wait for Clk_period;
		Addr <=  "0010010010010";
		Trees_din <= x"002c12ed";
		wait for Clk_period;
		Addr <=  "0010010010011";
		Trees_din <= x"cffff304";
		wait for Clk_period;
		Addr <=  "0010010010100";
		Trees_din <= x"008712ed";
		wait for Clk_period;
		Addr <=  "0010010010101";
		Trees_din <= x"ffaa12ed";
		wait for Clk_period;
		Addr <=  "0010010010110";
		Trees_din <= x"23ff2d08";
		wait for Clk_period;
		Addr <=  "0010010010111";
		Trees_din <= x"79fef104";
		wait for Clk_period;
		Addr <=  "0010010011000";
		Trees_din <= x"006712ed";
		wait for Clk_period;
		Addr <=  "0010010011001";
		Trees_din <= x"ffc212ed";
		wait for Clk_period;
		Addr <=  "0010010011010";
		Trees_din <= x"9c002e04";
		wait for Clk_period;
		Addr <=  "0010010011011";
		Trees_din <= x"ff7512ed";
		wait for Clk_period;
		Addr <=  "0010010011100";
		Trees_din <= x"fff612ed";
		wait for Clk_period;
		Addr <=  "0010010011101";
		Trees_din <= x"83ffbd10";
		wait for Clk_period;
		Addr <=  "0010010011110";
		Trees_din <= x"ee009c08";
		wait for Clk_period;
		Addr <=  "0010010011111";
		Trees_din <= x"7d004104";
		wait for Clk_period;
		Addr <=  "0010010100000";
		Trees_din <= x"ff6e12ed";
		wait for Clk_period;
		Addr <=  "0010010100001";
		Trees_din <= x"ffd412ed";
		wait for Clk_period;
		Addr <=  "0010010100010";
		Trees_din <= x"b5fea504";
		wait for Clk_period;
		Addr <=  "0010010100011";
		Trees_din <= x"006112ed";
		wait for Clk_period;
		Addr <=  "0010010100100";
		Trees_din <= x"ffad12ed";
		wait for Clk_period;
		Addr <=  "0010010100101";
		Trees_din <= x"5fff4008";
		wait for Clk_period;
		Addr <=  "0010010100110";
		Trees_din <= x"25005204";
		wait for Clk_period;
		Addr <=  "0010010100111";
		Trees_din <= x"fffb12ed";
		wait for Clk_period;
		Addr <=  "0010010101000";
		Trees_din <= x"00a412ed";
		wait for Clk_period;
		Addr <=  "0010010101001";
		Trees_din <= x"ffa612ed";
		wait for Clk_period;
		Addr <=  "0010010101010";
		Trees_din <= x"96ff3418";
		wait for Clk_period;
		Addr <=  "0010010101011";
		Trees_din <= x"fbff1c08";
		wait for Clk_period;
		Addr <=  "0010010101100";
		Trees_din <= x"24ffb104";
		wait for Clk_period;
		Addr <=  "0010010101101";
		Trees_din <= x"ffe712ed";
		wait for Clk_period;
		Addr <=  "0010010101110";
		Trees_din <= x"00a612ed";
		wait for Clk_period;
		Addr <=  "0010010101111";
		Trees_din <= x"53ffc504";
		wait for Clk_period;
		Addr <=  "0010010110000";
		Trees_din <= x"ff7d12ed";
		wait for Clk_period;
		Addr <=  "0010010110001";
		Trees_din <= x"9dff9a08";
		wait for Clk_period;
		Addr <=  "0010010110010";
		Trees_din <= x"bdfffe04";
		wait for Clk_period;
		Addr <=  "0010010110011";
		Trees_din <= x"ffec12ed";
		wait for Clk_period;
		Addr <=  "0010010110100";
		Trees_din <= x"009512ed";
		wait for Clk_period;
		Addr <=  "0010010110101";
		Trees_din <= x"ff9b12ed";
		wait for Clk_period;
		Addr <=  "0010010110110";
		Trees_din <= x"9ffe9504";
		wait for Clk_period;
		Addr <=  "0010010110111";
		Trees_din <= x"002212ed";
		wait for Clk_period;
		Addr <=  "0010010111000";
		Trees_din <= x"ef002404";
		wait for Clk_period;
		Addr <=  "0010010111001";
		Trees_din <= x"ff6b12ed";
		wait for Clk_period;
		Addr <=  "0010010111010";
		Trees_din <= x"000f12ed";
		wait for Clk_period;
		Addr <=  "0010010111011";
		Trees_din <= x"42ffa550";
		wait for Clk_period;
		Addr <=  "0010010111100";
		Trees_din <= x"c1fed328";
		wait for Clk_period;
		Addr <=  "0010010111101";
		Trees_din <= x"7500f01c";
		wait for Clk_period;
		Addr <=  "0010010111110";
		Trees_din <= x"8dfe6110";
		wait for Clk_period;
		Addr <=  "0010010111111";
		Trees_din <= x"2dfee508";
		wait for Clk_period;
		Addr <=  "0010011000000";
		Trees_din <= x"32fe8204";
		wait for Clk_period;
		Addr <=  "0010011000001";
		Trees_din <= x"ff8f13b9";
		wait for Clk_period;
		Addr <=  "0010011000010";
		Trees_din <= x"005c13b9";
		wait for Clk_period;
		Addr <=  "0010011000011";
		Trees_din <= x"4bfe1004";
		wait for Clk_period;
		Addr <=  "0010011000100";
		Trees_din <= x"002713b9";
		wait for Clk_period;
		Addr <=  "0010011000101";
		Trees_din <= x"ff7813b9";
		wait for Clk_period;
		Addr <=  "0010011000110";
		Trees_din <= x"31005504";
		wait for Clk_period;
		Addr <=  "0010011000111";
		Trees_din <= x"ff6d13b9";
		wait for Clk_period;
		Addr <=  "0010011001000";
		Trees_din <= x"26009804";
		wait for Clk_period;
		Addr <=  "0010011001001";
		Trees_din <= x"ffa113b9";
		wait for Clk_period;
		Addr <=  "0010011001010";
		Trees_din <= x"005d13b9";
		wait for Clk_period;
		Addr <=  "0010011001011";
		Trees_din <= x"52ff2004";
		wait for Clk_period;
		Addr <=  "0010011001100";
		Trees_din <= x"ffd813b9";
		wait for Clk_period;
		Addr <=  "0010011001101";
		Trees_din <= x"95ff2504";
		wait for Clk_period;
		Addr <=  "0010011001110";
		Trees_din <= x"003313b9";
		wait for Clk_period;
		Addr <=  "0010011001111";
		Trees_din <= x"00d113b9";
		wait for Clk_period;
		Addr <=  "0010011010000";
		Trees_din <= x"29ff7414";
		wait for Clk_period;
		Addr <=  "0010011010001";
		Trees_din <= x"51ff5108";
		wait for Clk_period;
		Addr <=  "0010011010010";
		Trees_din <= x"83ff5604";
		wait for Clk_period;
		Addr <=  "0010011010011";
		Trees_din <= x"ffa113b9";
		wait for Clk_period;
		Addr <=  "0010011010100";
		Trees_din <= x"ffe813b9";
		wait for Clk_period;
		Addr <=  "0010011010101";
		Trees_din <= x"64fedb04";
		wait for Clk_period;
		Addr <=  "0010011010110";
		Trees_din <= x"ffac13b9";
		wait for Clk_period;
		Addr <=  "0010011010111";
		Trees_din <= x"3f008204";
		wait for Clk_period;
		Addr <=  "0010011011000";
		Trees_din <= x"006f13b9";
		wait for Clk_period;
		Addr <=  "0010011011001";
		Trees_din <= x"ffbb13b9";
		wait for Clk_period;
		Addr <=  "0010011011010";
		Trees_din <= x"2900560c";
		wait for Clk_period;
		Addr <=  "0010011011011";
		Trees_din <= x"4afe7f04";
		wait for Clk_period;
		Addr <=  "0010011011100";
		Trees_din <= x"004d13b9";
		wait for Clk_period;
		Addr <=  "0010011011101";
		Trees_din <= x"06006304";
		wait for Clk_period;
		Addr <=  "0010011011110";
		Trees_din <= x"ff7413b9";
		wait for Clk_period;
		Addr <=  "0010011011111";
		Trees_din <= x"000a13b9";
		wait for Clk_period;
		Addr <=  "0010011100000";
		Trees_din <= x"d2feb904";
		wait for Clk_period;
		Addr <=  "0010011100001";
		Trees_din <= x"009513b9";
		wait for Clk_period;
		Addr <=  "0010011100010";
		Trees_din <= x"ffea13b9";
		wait for Clk_period;
		Addr <=  "0010011100011";
		Trees_din <= x"e2fea50c";
		wait for Clk_period;
		Addr <=  "0010011100100";
		Trees_din <= x"12ffe804";
		wait for Clk_period;
		Addr <=  "0010011100101";
		Trees_din <= x"ff9d13b9";
		wait for Clk_period;
		Addr <=  "0010011100110";
		Trees_din <= x"c0ff6804";
		wait for Clk_period;
		Addr <=  "0010011100111";
		Trees_din <= x"007d13b9";
		wait for Clk_period;
		Addr <=  "0010011101000";
		Trees_din <= x"ffdf13b9";
		wait for Clk_period;
		Addr <=  "0010011101001";
		Trees_din <= x"d2fe0304";
		wait for Clk_period;
		Addr <=  "0010011101010";
		Trees_din <= x"001e13b9";
		wait for Clk_period;
		Addr <=  "0010011101011";
		Trees_din <= x"4afe6a04";
		wait for Clk_period;
		Addr <=  "0010011101100";
		Trees_din <= x"001613b9";
		wait for Clk_period;
		Addr <=  "0010011101101";
		Trees_din <= x"ff6c13b9";
		wait for Clk_period;
		Addr <=  "0010011101110";
		Trees_din <= x"b8ff8640";
		wait for Clk_period;
		Addr <=  "0010011101111";
		Trees_din <= x"b4ff1a24";
		wait for Clk_period;
		Addr <=  "0010011110000";
		Trees_din <= x"78ffd41c";
		wait for Clk_period;
		Addr <=  "0010011110001";
		Trees_din <= x"58fed010";
		wait for Clk_period;
		Addr <=  "0010011110010";
		Trees_din <= x"faffb808";
		wait for Clk_period;
		Addr <=  "0010011110011";
		Trees_din <= x"68ff9e04";
		wait for Clk_period;
		Addr <=  "0010011110100";
		Trees_din <= x"ff7e147d";
		wait for Clk_period;
		Addr <=  "0010011110101";
		Trees_din <= x"003b147d";
		wait for Clk_period;
		Addr <=  "0010011110110";
		Trees_din <= x"adff4c04";
		wait for Clk_period;
		Addr <=  "0010011110111";
		Trees_din <= x"008f147d";
		wait for Clk_period;
		Addr <=  "0010011111000";
		Trees_din <= x"ffb9147d";
		wait for Clk_period;
		Addr <=  "0010011111001";
		Trees_din <= x"b3ff7908";
		wait for Clk_period;
		Addr <=  "0010011111010";
		Trees_din <= x"a4ff7204";
		wait for Clk_period;
		Addr <=  "0010011111011";
		Trees_din <= x"ffff147d";
		wait for Clk_period;
		Addr <=  "0010011111100";
		Trees_din <= x"0067147d";
		wait for Clk_period;
		Addr <=  "0010011111101";
		Trees_din <= x"ff98147d";
		wait for Clk_period;
		Addr <=  "0010011111110";
		Trees_din <= x"5fffa604";
		wait for Clk_period;
		Addr <=  "0010011111111";
		Trees_din <= x"ff7f147d";
		wait for Clk_period;
		Addr <=  "0010100000000";
		Trees_din <= x"ffea147d";
		wait for Clk_period;
		Addr <=  "0010100000001";
		Trees_din <= x"83ffbd10";
		wait for Clk_period;
		Addr <=  "0010100000010";
		Trees_din <= x"ee009c08";
		wait for Clk_period;
		Addr <=  "0010100000011";
		Trees_din <= x"43fee704";
		wait for Clk_period;
		Addr <=  "0010100000100";
		Trees_din <= x"ffdf147d";
		wait for Clk_period;
		Addr <=  "0010100000101";
		Trees_din <= x"ff71147d";
		wait for Clk_period;
		Addr <=  "0010100000110";
		Trees_din <= x"52fecf04";
		wait for Clk_period;
		Addr <=  "0010100000111";
		Trees_din <= x"0058147d";
		wait for Clk_period;
		Addr <=  "0010100001000";
		Trees_din <= x"ffd0147d";
		wait for Clk_period;
		Addr <=  "0010100001001";
		Trees_din <= x"5fff4008";
		wait for Clk_period;
		Addr <=  "0010100001010";
		Trees_din <= x"75003904";
		wait for Clk_period;
		Addr <=  "0010100001011";
		Trees_din <= x"000d147d";
		wait for Clk_period;
		Addr <=  "0010100001100";
		Trees_din <= x"0090147d";
		wait for Clk_period;
		Addr <=  "0010100001101";
		Trees_din <= x"ffaf147d";
		wait for Clk_period;
		Addr <=  "0010100001110";
		Trees_din <= x"96ff3418";
		wait for Clk_period;
		Addr <=  "0010100001111";
		Trees_din <= x"fbff0d08";
		wait for Clk_period;
		Addr <=  "0010100010000";
		Trees_din <= x"b5ff1504";
		wait for Clk_period;
		Addr <=  "0010100010001";
		Trees_din <= x"0007147d";
		wait for Clk_period;
		Addr <=  "0010100010010";
		Trees_din <= x"009a147d";
		wait for Clk_period;
		Addr <=  "0010100010011";
		Trees_din <= x"cafef50c";
		wait for Clk_period;
		Addr <=  "0010100010100";
		Trees_din <= x"f5ff6c04";
		wait for Clk_period;
		Addr <=  "0010100010101";
		Trees_din <= x"0049147d";
		wait for Clk_period;
		Addr <=  "0010100010110";
		Trees_din <= x"a4ff1b04";
		wait for Clk_period;
		Addr <=  "0010100010111";
		Trees_din <= x"0008147d";
		wait for Clk_period;
		Addr <=  "0010100011000";
		Trees_din <= x"ff78147d";
		wait for Clk_period;
		Addr <=  "0010100011001";
		Trees_din <= x"0065147d";
		wait for Clk_period;
		Addr <=  "0010100011010";
		Trees_din <= x"30003604";
		wait for Clk_period;
		Addr <=  "0010100011011";
		Trees_din <= x"ff6e147d";
		wait for Clk_period;
		Addr <=  "0010100011100";
		Trees_din <= x"03000104";
		wait for Clk_period;
		Addr <=  "0010100011101";
		Trees_din <= x"ff98147d";
		wait for Clk_period;
		Addr <=  "0010100011110";
		Trees_din <= x"0056147d";
		wait for Clk_period;
		Addr <=  "0010100011111";
		Trees_din <= x"42ffa53c";
		wait for Clk_period;
		Addr <=  "0010100100000";
		Trees_din <= x"58fea914";
		wait for Clk_period;
		Addr <=  "0010100100001";
		Trees_din <= x"1aff1b08";
		wait for Clk_period;
		Addr <=  "0010100100010";
		Trees_din <= x"c2fed204";
		wait for Clk_period;
		Addr <=  "0010100100011";
		Trees_din <= x"fff71521";
		wait for Clk_period;
		Addr <=  "0010100100100";
		Trees_din <= x"ff751521";
		wait for Clk_period;
		Addr <=  "0010100100101";
		Trees_din <= x"77fecb08";
		wait for Clk_period;
		Addr <=  "0010100100110";
		Trees_din <= x"56ff5f04";
		wait for Clk_period;
		Addr <=  "0010100100111";
		Trees_din <= x"00891521";
		wait for Clk_period;
		Addr <=  "0010100101000";
		Trees_din <= x"ffd81521";
		wait for Clk_period;
		Addr <=  "0010100101001";
		Trees_din <= x"ff9a1521";
		wait for Clk_period;
		Addr <=  "0010100101010";
		Trees_din <= x"75ffaf08";
		wait for Clk_period;
		Addr <=  "0010100101011";
		Trees_din <= x"51005004";
		wait for Clk_period;
		Addr <=  "0010100101100";
		Trees_din <= x"ff801521";
		wait for Clk_period;
		Addr <=  "0010100101101";
		Trees_din <= x"00021521";
		wait for Clk_period;
		Addr <=  "0010100101110";
		Trees_din <= x"79ff1310";
		wait for Clk_period;
		Addr <=  "0010100101111";
		Trees_din <= x"46feaf08";
		wait for Clk_period;
		Addr <=  "0010100110000";
		Trees_din <= x"cd002e04";
		wait for Clk_period;
		Addr <=  "0010100110001";
		Trees_din <= x"ff991521";
		wait for Clk_period;
		Addr <=  "0010100110010";
		Trees_din <= x"00121521";
		wait for Clk_period;
		Addr <=  "0010100110011";
		Trees_din <= x"eeff9c04";
		wait for Clk_period;
		Addr <=  "0010100110100";
		Trees_din <= x"ffc71521";
		wait for Clk_period;
		Addr <=  "0010100110101";
		Trees_din <= x"00731521";
		wait for Clk_period;
		Addr <=  "0010100110110";
		Trees_din <= x"adff9e08";
		wait for Clk_period;
		Addr <=  "0010100110111";
		Trees_din <= x"25009104";
		wait for Clk_period;
		Addr <=  "0010100111000";
		Trees_din <= x"ffec1521";
		wait for Clk_period;
		Addr <=  "0010100111001";
		Trees_din <= x"005e1521";
		wait for Clk_period;
		Addr <=  "0010100111010";
		Trees_din <= x"eeff4004";
		wait for Clk_period;
		Addr <=  "0010100111011";
		Trees_din <= x"00301521";
		wait for Clk_period;
		Addr <=  "0010100111100";
		Trees_din <= x"ff7e1521";
		wait for Clk_period;
		Addr <=  "0010100111101";
		Trees_din <= x"14fe4c08";
		wait for Clk_period;
		Addr <=  "0010100111110";
		Trees_din <= x"aefe7104";
		wait for Clk_period;
		Addr <=  "0010100111111";
		Trees_din <= x"00691521";
		wait for Clk_period;
		Addr <=  "0010101000000";
		Trees_din <= x"ffcc1521";
		wait for Clk_period;
		Addr <=  "0010101000001";
		Trees_din <= x"dc005008";
		wait for Clk_period;
		Addr <=  "0010101000010";
		Trees_din <= x"1f00df04";
		wait for Clk_period;
		Addr <=  "0010101000011";
		Trees_din <= x"ff6f1521";
		wait for Clk_period;
		Addr <=  "0010101000100";
		Trees_din <= x"ffe61521";
		wait for Clk_period;
		Addr <=  "0010101000101";
		Trees_din <= x"ebfe9a04";
		wait for Clk_period;
		Addr <=  "0010101000110";
		Trees_din <= x"00451521";
		wait for Clk_period;
		Addr <=  "0010101000111";
		Trees_din <= x"ffa71521";
		wait for Clk_period;
		Addr <=  "0010101001000";
		Trees_din <= x"9eff7828";
		wait for Clk_period;
		Addr <=  "0010101001001";
		Trees_din <= x"6bff1320";
		wait for Clk_period;
		Addr <=  "0010101001010";
		Trees_din <= x"c0ffa818";
		wait for Clk_period;
		Addr <=  "0010101001011";
		Trees_din <= x"c0ff180c";
		wait for Clk_period;
		Addr <=  "0010101001100";
		Trees_din <= x"15001f08";
		wait for Clk_period;
		Addr <=  "0010101001101";
		Trees_din <= x"b0ffb504";
		wait for Clk_period;
		Addr <=  "0010101001110";
		Trees_din <= x"ff8115bd";
		wait for Clk_period;
		Addr <=  "0010101001111";
		Trees_din <= x"000515bd";
		wait for Clk_period;
		Addr <=  "0010101010000";
		Trees_din <= x"004415bd";
		wait for Clk_period;
		Addr <=  "0010101010001";
		Trees_din <= x"76ff5104";
		wait for Clk_period;
		Addr <=  "0010101010010";
		Trees_din <= x"ff9415bd";
		wait for Clk_period;
		Addr <=  "0010101010011";
		Trees_din <= x"adffa404";
		wait for Clk_period;
		Addr <=  "0010101010100";
		Trees_din <= x"005315bd";
		wait for Clk_period;
		Addr <=  "0010101010101";
		Trees_din <= x"ffe815bd";
		wait for Clk_period;
		Addr <=  "0010101010110";
		Trees_din <= x"74ff8404";
		wait for Clk_period;
		Addr <=  "0010101010111";
		Trees_din <= x"001715bd";
		wait for Clk_period;
		Addr <=  "0010101011000";
		Trees_din <= x"ff8515bd";
		wait for Clk_period;
		Addr <=  "0010101011001";
		Trees_din <= x"57fe6b04";
		wait for Clk_period;
		Addr <=  "0010101011010";
		Trees_din <= x"002f15bd";
		wait for Clk_period;
		Addr <=  "0010101011011";
		Trees_din <= x"ff7a15bd";
		wait for Clk_period;
		Addr <=  "0010101011100";
		Trees_din <= x"23ff9e24";
		wait for Clk_period;
		Addr <=  "0010101011101";
		Trees_din <= x"baff620c";
		wait for Clk_period;
		Addr <=  "0010101011110";
		Trees_din <= x"0cfe8408";
		wait for Clk_period;
		Addr <=  "0010101011111";
		Trees_din <= x"00ff6e04";
		wait for Clk_period;
		Addr <=  "0010101100000";
		Trees_din <= x"000f15bd";
		wait for Clk_period;
		Addr <=  "0010101100001";
		Trees_din <= x"009d15bd";
		wait for Clk_period;
		Addr <=  "0010101100010";
		Trees_din <= x"ffaa15bd";
		wait for Clk_period;
		Addr <=  "0010101100011";
		Trees_din <= x"1cffbc08";
		wait for Clk_period;
		Addr <=  "0010101100100";
		Trees_din <= x"d2fe3304";
		wait for Clk_period;
		Addr <=  "0010101100101";
		Trees_din <= x"000d15bd";
		wait for Clk_period;
		Addr <=  "0010101100110";
		Trees_din <= x"ff7415bd";
		wait for Clk_period;
		Addr <=  "0010101100111";
		Trees_din <= x"b7ff5908";
		wait for Clk_period;
		Addr <=  "0010101101000";
		Trees_din <= x"60ff5404";
		wait for Clk_period;
		Addr <=  "0010101101001";
		Trees_din <= x"007715bd";
		wait for Clk_period;
		Addr <=  "0010101101010";
		Trees_din <= x"001915bd";
		wait for Clk_period;
		Addr <=  "0010101101011";
		Trees_din <= x"ceff8a04";
		wait for Clk_period;
		Addr <=  "0010101101100";
		Trees_din <= x"000f15bd";
		wait for Clk_period;
		Addr <=  "0010101101101";
		Trees_din <= x"ffaa15bd";
		wait for Clk_period;
		Addr <=  "0010101101110";
		Trees_din <= x"ff7515bd";
		wait for Clk_period;
		Addr <=  "0010101101111";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0010101110000";
		Trees_din <= x"42ffa548";
		wait for Clk_period;
		Addr <=  "0010101110001";
		Trees_din <= x"c1fed530";
		wait for Clk_period;
		Addr <=  "0010101110010";
		Trees_din <= x"66004920";
		wait for Clk_period;
		Addr <=  "0010101110011";
		Trees_din <= x"2fff1110";
		wait for Clk_period;
		Addr <=  "0010101110100";
		Trees_din <= x"80fff008";
		wait for Clk_period;
		Addr <=  "0010101110101";
		Trees_din <= x"65ffc104";
		wait for Clk_period;
		Addr <=  "0010101110110";
		Trees_din <= x"ff96167d";
		wait for Clk_period;
		Addr <=  "0010101110111";
		Trees_din <= x"003f167d";
		wait for Clk_period;
		Addr <=  "0010101111000";
		Trees_din <= x"59ff5104";
		wait for Clk_period;
		Addr <=  "0010101111001";
		Trees_din <= x"008e167d";
		wait for Clk_period;
		Addr <=  "0010101111010";
		Trees_din <= x"001a167d";
		wait for Clk_period;
		Addr <=  "0010101111011";
		Trees_din <= x"ce002708";
		wait for Clk_period;
		Addr <=  "0010101111100";
		Trees_din <= x"01fdf704";
		wait for Clk_period;
		Addr <=  "0010101111101";
		Trees_din <= x"0003167d";
		wait for Clk_period;
		Addr <=  "0010101111110";
		Trees_din <= x"ff76167d";
		wait for Clk_period;
		Addr <=  "0010101111111";
		Trees_din <= x"33ffcc04";
		wait for Clk_period;
		Addr <=  "0010110000000";
		Trees_din <= x"ffb9167d";
		wait for Clk_period;
		Addr <=  "0010110000001";
		Trees_din <= x"005f167d";
		wait for Clk_period;
		Addr <=  "0010110000010";
		Trees_din <= x"58fef708";
		wait for Clk_period;
		Addr <=  "0010110000011";
		Trees_din <= x"4afea804";
		wait for Clk_period;
		Addr <=  "0010110000100";
		Trees_din <= x"000c167d";
		wait for Clk_period;
		Addr <=  "0010110000101";
		Trees_din <= x"ffa2167d";
		wait for Clk_period;
		Addr <=  "0010110000110";
		Trees_din <= x"5dffe304";
		wait for Clk_period;
		Addr <=  "0010110000111";
		Trees_din <= x"009d167d";
		wait for Clk_period;
		Addr <=  "0010110001000";
		Trees_din <= x"fffb167d";
		wait for Clk_period;
		Addr <=  "0010110001001";
		Trees_din <= x"38ffd110";
		wait for Clk_period;
		Addr <=  "0010110001010";
		Trees_din <= x"64fedb04";
		wait for Clk_period;
		Addr <=  "0010110001011";
		Trees_din <= x"ffae167d";
		wait for Clk_period;
		Addr <=  "0010110001100";
		Trees_din <= x"3cff5e08";
		wait for Clk_period;
		Addr <=  "0010110001101";
		Trees_din <= x"98feb504";
		wait for Clk_period;
		Addr <=  "0010110001110";
		Trees_din <= x"ffff167d";
		wait for Clk_period;
		Addr <=  "0010110001111";
		Trees_din <= x"006e167d";
		wait for Clk_period;
		Addr <=  "0010110010000";
		Trees_din <= x"ffb4167d";
		wait for Clk_period;
		Addr <=  "0010110010001";
		Trees_din <= x"11fefc04";
		wait for Clk_period;
		Addr <=  "0010110010010";
		Trees_din <= x"002e167d";
		wait for Clk_period;
		Addr <=  "0010110010011";
		Trees_din <= x"ff90167d";
		wait for Clk_period;
		Addr <=  "0010110010100";
		Trees_din <= x"e2fec00c";
		wait for Clk_period;
		Addr <=  "0010110010101";
		Trees_din <= x"adff7f08";
		wait for Clk_period;
		Addr <=  "0010110010110";
		Trees_din <= x"aefe9f04";
		wait for Clk_period;
		Addr <=  "0010110010111";
		Trees_din <= x"0069167d";
		wait for Clk_period;
		Addr <=  "0010110011000";
		Trees_din <= x"ffd9167d";
		wait for Clk_period;
		Addr <=  "0010110011001";
		Trees_din <= x"ffa4167d";
		wait for Clk_period;
		Addr <=  "0010110011010";
		Trees_din <= x"d2fe0304";
		wait for Clk_period;
		Addr <=  "0010110011011";
		Trees_din <= x"0015167d";
		wait for Clk_period;
		Addr <=  "0010110011100";
		Trees_din <= x"c5ffbe04";
		wait for Clk_period;
		Addr <=  "0010110011101";
		Trees_din <= x"ff71167d";
		wait for Clk_period;
		Addr <=  "0010110011110";
		Trees_din <= x"ffe5167d";
		wait for Clk_period;
		Addr <=  "0010110011111";
		Trees_din <= x"29ff7948";
		wait for Clk_period;
		Addr <=  "0010110100000";
		Trees_din <= x"c1fed328";
		wait for Clk_period;
		Addr <=  "0010110100001";
		Trees_din <= x"66002b18";
		wait for Clk_period;
		Addr <=  "0010110100010";
		Trees_din <= x"80fffd10";
		wait for Clk_period;
		Addr <=  "0010110100011";
		Trees_din <= x"cdff6108";
		wait for Clk_period;
		Addr <=  "0010110100100";
		Trees_din <= x"63ff3f04";
		wait for Clk_period;
		Addr <=  "0010110100101";
		Trees_din <= x"004d1749";
		wait for Clk_period;
		Addr <=  "0010110100110";
		Trees_din <= x"ffb21749";
		wait for Clk_period;
		Addr <=  "0010110100111";
		Trees_din <= x"f5ff7d04";
		wait for Clk_period;
		Addr <=  "0010110101000";
		Trees_din <= x"000d1749";
		wait for Clk_period;
		Addr <=  "0010110101001";
		Trees_din <= x"ff721749";
		wait for Clk_period;
		Addr <=  "0010110101010";
		Trees_din <= x"8dfde004";
		wait for Clk_period;
		Addr <=  "0010110101011";
		Trees_din <= x"00821749";
		wait for Clk_period;
		Addr <=  "0010110101100";
		Trees_din <= x"ffd91749";
		wait for Clk_period;
		Addr <=  "0010110101101";
		Trees_din <= x"73ffde04";
		wait for Clk_period;
		Addr <=  "0010110101110";
		Trees_din <= x"ffcd1749";
		wait for Clk_period;
		Addr <=  "0010110101111";
		Trees_din <= x"ec000708";
		wait for Clk_period;
		Addr <=  "0010110110000";
		Trees_din <= x"eefff004";
		wait for Clk_period;
		Addr <=  "0010110110001";
		Trees_din <= x"001f1749";
		wait for Clk_period;
		Addr <=  "0010110110010";
		Trees_din <= x"008f1749";
		wait for Clk_period;
		Addr <=  "0010110110011";
		Trees_din <= x"ffee1749";
		wait for Clk_period;
		Addr <=  "0010110110100";
		Trees_din <= x"16ff3e10";
		wait for Clk_period;
		Addr <=  "0010110110101";
		Trees_din <= x"b8ffbf0c";
		wait for Clk_period;
		Addr <=  "0010110110110";
		Trees_din <= x"dfffe608";
		wait for Clk_period;
		Addr <=  "0010110110111";
		Trees_din <= x"fb001204";
		wait for Clk_period;
		Addr <=  "0010110111000";
		Trees_din <= x"00691749";
		wait for Clk_period;
		Addr <=  "0010110111001";
		Trees_din <= x"ffd91749";
		wait for Clk_period;
		Addr <=  "0010110111010";
		Trees_din <= x"ffb21749";
		wait for Clk_period;
		Addr <=  "0010110111011";
		Trees_din <= x"ffa31749";
		wait for Clk_period;
		Addr <=  "0010110111100";
		Trees_din <= x"f7ff0408";
		wait for Clk_period;
		Addr <=  "0010110111101";
		Trees_din <= x"84ffdc04";
		wait for Clk_period;
		Addr <=  "0010110111110";
		Trees_din <= x"ffed1749";
		wait for Clk_period;
		Addr <=  "0010110111111";
		Trees_din <= x"004c1749";
		wait for Clk_period;
		Addr <=  "0010111000000";
		Trees_din <= x"6aff3f04";
		wait for Clk_period;
		Addr <=  "0010111000001";
		Trees_din <= x"ffea1749";
		wait for Clk_period;
		Addr <=  "0010111000010";
		Trees_din <= x"ff8e1749";
		wait for Clk_period;
		Addr <=  "0010111000011";
		Trees_din <= x"2700050c";
		wait for Clk_period;
		Addr <=  "0010111000100";
		Trees_din <= x"ec006a08";
		wait for Clk_period;
		Addr <=  "0010111000101";
		Trees_din <= x"81fef504";
		wait for Clk_period;
		Addr <=  "0010111000110";
		Trees_din <= x"ffea1749";
		wait for Clk_period;
		Addr <=  "0010111000111";
		Trees_din <= x"ff711749";
		wait for Clk_period;
		Addr <=  "0010111001000";
		Trees_din <= x"001c1749";
		wait for Clk_period;
		Addr <=  "0010111001001";
		Trees_din <= x"adff8310";
		wait for Clk_period;
		Addr <=  "0010111001010";
		Trees_din <= x"8effd104";
		wait for Clk_period;
		Addr <=  "0010111001011";
		Trees_din <= x"ffa91749";
		wait for Clk_period;
		Addr <=  "0010111001100";
		Trees_din <= x"68febd04";
		wait for Clk_period;
		Addr <=  "0010111001101";
		Trees_din <= x"ffc41749";
		wait for Clk_period;
		Addr <=  "0010111001110";
		Trees_din <= x"46fee904";
		wait for Clk_period;
		Addr <=  "0010111001111";
		Trees_din <= x"fff11749";
		wait for Clk_period;
		Addr <=  "0010111010000";
		Trees_din <= x"007d1749";
		wait for Clk_period;
		Addr <=  "0010111010001";
		Trees_din <= x"ff8c1749";
		wait for Clk_period;
		Addr <=  "0010111010010";
		Trees_din <= x"29ff7948";
		wait for Clk_period;
		Addr <=  "0010111010011";
		Trees_din <= x"8dfe0f1c";
		wait for Clk_period;
		Addr <=  "0010111010100";
		Trees_din <= x"58fed50c";
		wait for Clk_period;
		Addr <=  "0010111010101";
		Trees_din <= x"55000708";
		wait for Clk_period;
		Addr <=  "0010111010110";
		Trees_din <= x"b7ff0904";
		wait for Clk_period;
		Addr <=  "0010111010111";
		Trees_din <= x"0055181d";
		wait for Clk_period;
		Addr <=  "0010111011000";
		Trees_din <= x"fff0181d";
		wait for Clk_period;
		Addr <=  "0010111011001";
		Trees_din <= x"ff95181d";
		wait for Clk_period;
		Addr <=  "0010111011010";
		Trees_din <= x"7a00050c";
		wait for Clk_period;
		Addr <=  "0010111011011";
		Trees_din <= x"a3ff8e08";
		wait for Clk_period;
		Addr <=  "0010111011100";
		Trees_din <= x"aeff2904";
		wait for Clk_period;
		Addr <=  "0010111011101";
		Trees_din <= x"0088181d";
		wait for Clk_period;
		Addr <=  "0010111011110";
		Trees_din <= x"0014181d";
		wait for Clk_period;
		Addr <=  "0010111011111";
		Trees_din <= x"fff6181d";
		wait for Clk_period;
		Addr <=  "0010111100000";
		Trees_din <= x"ffcc181d";
		wait for Clk_period;
		Addr <=  "0010111100001";
		Trees_din <= x"aeff2f18";
		wait for Clk_period;
		Addr <=  "0010111100010";
		Trees_din <= x"25002908";
		wait for Clk_period;
		Addr <=  "0010111100011";
		Trees_din <= x"b5ff5304";
		wait for Clk_period;
		Addr <=  "0010111100100";
		Trees_din <= x"ff78181d";
		wait for Clk_period;
		Addr <=  "0010111100101";
		Trees_din <= x"ffeb181d";
		wait for Clk_period;
		Addr <=  "0010111100110";
		Trees_din <= x"98ff3308";
		wait for Clk_period;
		Addr <=  "0010111100111";
		Trees_din <= x"e2fefb04";
		wait for Clk_period;
		Addr <=  "0010111101000";
		Trees_din <= x"0007181d";
		wait for Clk_period;
		Addr <=  "0010111101001";
		Trees_din <= x"ff92181d";
		wait for Clk_period;
		Addr <=  "0010111101010";
		Trees_din <= x"a2ff9204";
		wait for Clk_period;
		Addr <=  "0010111101011";
		Trees_din <= x"006b181d";
		wait for Clk_period;
		Addr <=  "0010111101100";
		Trees_din <= x"fff7181d";
		wait for Clk_period;
		Addr <=  "0010111101101";
		Trees_din <= x"b1ff0f0c";
		wait for Clk_period;
		Addr <=  "0010111101110";
		Trees_din <= x"18ff8204";
		wait for Clk_period;
		Addr <=  "0010111101111";
		Trees_din <= x"ffc1181d";
		wait for Clk_period;
		Addr <=  "0010111110000";
		Trees_din <= x"f6fedb04";
		wait for Clk_period;
		Addr <=  "0010111110001";
		Trees_din <= x"0001181d";
		wait for Clk_period;
		Addr <=  "0010111110010";
		Trees_din <= x"0097181d";
		wait for Clk_period;
		Addr <=  "0010111110011";
		Trees_din <= x"66004404";
		wait for Clk_period;
		Addr <=  "0010111110100";
		Trees_din <= x"ff8b181d";
		wait for Clk_period;
		Addr <=  "0010111110101";
		Trees_din <= x"0038181d";
		wait for Clk_period;
		Addr <=  "0010111110110";
		Trees_din <= x"2900561c";
		wait for Clk_period;
		Addr <=  "0010111110111";
		Trees_din <= x"4afe7f08";
		wait for Clk_period;
		Addr <=  "0010111111000";
		Trees_din <= x"e8ff7b04";
		wait for Clk_period;
		Addr <=  "0010111111001";
		Trees_din <= x"005e181d";
		wait for Clk_period;
		Addr <=  "0010111111010";
		Trees_din <= x"ffb0181d";
		wait for Clk_period;
		Addr <=  "0010111111011";
		Trees_din <= x"b1fe9208";
		wait for Clk_period;
		Addr <=  "0010111111100";
		Trees_din <= x"18005304";
		wait for Clk_period;
		Addr <=  "0010111111101";
		Trees_din <= x"ffa6181d";
		wait for Clk_period;
		Addr <=  "0010111111110";
		Trees_din <= x"0050181d";
		wait for Clk_period;
		Addr <=  "0010111111111";
		Trees_din <= x"3b000008";
		wait for Clk_period;
		Addr <=  "0011000000000";
		Trees_din <= x"1bff0f04";
		wait for Clk_period;
		Addr <=  "0011000000001";
		Trees_din <= x"ffe1181d";
		wait for Clk_period;
		Addr <=  "0011000000010";
		Trees_din <= x"ff70181d";
		wait for Clk_period;
		Addr <=  "0011000000011";
		Trees_din <= x"0009181d";
		wait for Clk_period;
		Addr <=  "0011000000100";
		Trees_din <= x"1f001504";
		wait for Clk_period;
		Addr <=  "0011000000101";
		Trees_din <= x"ffd5181d";
		wait for Clk_period;
		Addr <=  "0011000000110";
		Trees_din <= x"0077181d";
		wait for Clk_period;
		Addr <=  "0011000000111";
		Trees_din <= x"27000538";
		wait for Clk_period;
		Addr <=  "0011000001000";
		Trees_din <= x"29ff792c";
		wait for Clk_period;
		Addr <=  "0011000001001";
		Trees_din <= x"98feeb14";
		wait for Clk_period;
		Addr <=  "0011000001010";
		Trees_din <= x"6afff708";
		wait for Clk_period;
		Addr <=  "0011000001011";
		Trees_din <= x"0b009904";
		wait for Clk_period;
		Addr <=  "0011000001100";
		Trees_din <= x"ff7d18f1";
		wait for Clk_period;
		Addr <=  "0011000001101";
		Trees_din <= x"001718f1";
		wait for Clk_period;
		Addr <=  "0011000001110";
		Trees_din <= x"bdff1104";
		wait for Clk_period;
		Addr <=  "0011000001111";
		Trees_din <= x"007618f1";
		wait for Clk_period;
		Addr <=  "0011000010000";
		Trees_din <= x"47005204";
		wait for Clk_period;
		Addr <=  "0011000010001";
		Trees_din <= x"ffca18f1";
		wait for Clk_period;
		Addr <=  "0011000010010";
		Trees_din <= x"001a18f1";
		wait for Clk_period;
		Addr <=  "0011000010011";
		Trees_din <= x"45fee408";
		wait for Clk_period;
		Addr <=  "0011000010100";
		Trees_din <= x"0500ab04";
		wait for Clk_period;
		Addr <=  "0011000010101";
		Trees_din <= x"ff9118f1";
		wait for Clk_period;
		Addr <=  "0011000010110";
		Trees_din <= x"002c18f1";
		wait for Clk_period;
		Addr <=  "0011000010111";
		Trees_din <= x"13010908";
		wait for Clk_period;
		Addr <=  "0011000011000";
		Trees_din <= x"c1fee304";
		wait for Clk_period;
		Addr <=  "0011000011001";
		Trees_din <= x"001518f1";
		wait for Clk_period;
		Addr <=  "0011000011010";
		Trees_din <= x"008918f1";
		wait for Clk_period;
		Addr <=  "0011000011011";
		Trees_din <= x"e7ffe204";
		wait for Clk_period;
		Addr <=  "0011000011100";
		Trees_din <= x"ffab18f1";
		wait for Clk_period;
		Addr <=  "0011000011101";
		Trees_din <= x"003518f1";
		wait for Clk_period;
		Addr <=  "0011000011110";
		Trees_din <= x"6c000304";
		wait for Clk_period;
		Addr <=  "0011000011111";
		Trees_din <= x"ff7518f1";
		wait for Clk_period;
		Addr <=  "0011000100000";
		Trees_din <= x"46ff5604";
		wait for Clk_period;
		Addr <=  "0011000100001";
		Trees_din <= x"ffb218f1";
		wait for Clk_period;
		Addr <=  "0011000100010";
		Trees_din <= x"004d18f1";
		wait for Clk_period;
		Addr <=  "0011000100011";
		Trees_din <= x"15ffa114";
		wait for Clk_period;
		Addr <=  "0011000100100";
		Trees_din <= x"c0ff5e08";
		wait for Clk_period;
		Addr <=  "0011000100101";
		Trees_din <= x"e6ff5904";
		wait for Clk_period;
		Addr <=  "0011000100110";
		Trees_din <= x"000918f1";
		wait for Clk_period;
		Addr <=  "0011000100111";
		Trees_din <= x"ff8218f1";
		wait for Clk_period;
		Addr <=  "0011000101000";
		Trees_din <= x"f4fed008";
		wait for Clk_period;
		Addr <=  "0011000101001";
		Trees_din <= x"92ff2104";
		wait for Clk_period;
		Addr <=  "0011000101010";
		Trees_din <= x"000118f1";
		wait for Clk_period;
		Addr <=  "0011000101011";
		Trees_din <= x"007818f1";
		wait for Clk_period;
		Addr <=  "0011000101100";
		Trees_din <= x"ffa118f1";
		wait for Clk_period;
		Addr <=  "0011000101101";
		Trees_din <= x"32fe8208";
		wait for Clk_period;
		Addr <=  "0011000101110";
		Trees_din <= x"2a00c604";
		wait for Clk_period;
		Addr <=  "0011000101111";
		Trees_din <= x"ffa818f1";
		wait for Clk_period;
		Addr <=  "0011000110000";
		Trees_din <= x"002e18f1";
		wait for Clk_period;
		Addr <=  "0011000110001";
		Trees_din <= x"2dfee20c";
		wait for Clk_period;
		Addr <=  "0011000110010";
		Trees_din <= x"d1ff2004";
		wait for Clk_period;
		Addr <=  "0011000110011";
		Trees_din <= x"ffee18f1";
		wait for Clk_period;
		Addr <=  "0011000110100";
		Trees_din <= x"21ffd204";
		wait for Clk_period;
		Addr <=  "0011000110101";
		Trees_din <= x"008518f1";
		wait for Clk_period;
		Addr <=  "0011000110110";
		Trees_din <= x"000018f1";
		wait for Clk_period;
		Addr <=  "0011000110111";
		Trees_din <= x"e2fee908";
		wait for Clk_period;
		Addr <=  "0011000111000";
		Trees_din <= x"6d006004";
		wait for Clk_period;
		Addr <=  "0011000111001";
		Trees_din <= x"ffe718f1";
		wait for Clk_period;
		Addr <=  "0011000111010";
		Trees_din <= x"005d18f1";
		wait for Clk_period;
		Addr <=  "0011000111011";
		Trees_din <= x"ffa918f1";
		wait for Clk_period;
		Addr <=  "0011000111100";
		Trees_din <= x"25001920";
		wait for Clk_period;
		Addr <=  "0011000111101";
		Trees_din <= x"28feaf0c";
		wait for Clk_period;
		Addr <=  "0011000111110";
		Trees_din <= x"80ff9904";
		wait for Clk_period;
		Addr <=  "0011000111111";
		Trees_din <= x"ffa41995";
		wait for Clk_period;
		Addr <=  "0011001000000";
		Trees_din <= x"35fe9204";
		wait for Clk_period;
		Addr <=  "0011001000001";
		Trees_din <= x"00781995";
		wait for Clk_period;
		Addr <=  "0011001000010";
		Trees_din <= x"00111995";
		wait for Clk_period;
		Addr <=  "0011001000011";
		Trees_din <= x"68fe2f08";
		wait for Clk_period;
		Addr <=  "0011001000100";
		Trees_din <= x"ecff3f04";
		wait for Clk_period;
		Addr <=  "0011001000101";
		Trees_din <= x"00841995";
		wait for Clk_period;
		Addr <=  "0011001000110";
		Trees_din <= x"ffd51995";
		wait for Clk_period;
		Addr <=  "0011001000111";
		Trees_din <= x"b7fedc04";
		wait for Clk_period;
		Addr <=  "0011001001000";
		Trees_din <= x"00241995";
		wait for Clk_period;
		Addr <=  "0011001001001";
		Trees_din <= x"0b006504";
		wait for Clk_period;
		Addr <=  "0011001001010";
		Trees_din <= x"ff711995";
		wait for Clk_period;
		Addr <=  "0011001001011";
		Trees_din <= x"ffdf1995";
		wait for Clk_period;
		Addr <=  "0011001001100";
		Trees_din <= x"4aff4928";
		wait for Clk_period;
		Addr <=  "0011001001101";
		Trees_din <= x"2dff3418";
		wait for Clk_period;
		Addr <=  "0011001001110";
		Trees_din <= x"46fec908";
		wait for Clk_period;
		Addr <=  "0011001001111";
		Trees_din <= x"21000104";
		wait for Clk_period;
		Addr <=  "0011001010000";
		Trees_din <= x"ff961995";
		wait for Clk_period;
		Addr <=  "0011001010001";
		Trees_din <= x"00451995";
		wait for Clk_period;
		Addr <=  "0011001010010";
		Trees_din <= x"8aff8308";
		wait for Clk_period;
		Addr <=  "0011001010011";
		Trees_din <= x"16ff3304";
		wait for Clk_period;
		Addr <=  "0011001010100";
		Trees_din <= x"ffb21995";
		wait for Clk_period;
		Addr <=  "0011001010101";
		Trees_din <= x"003e1995";
		wait for Clk_period;
		Addr <=  "0011001010110";
		Trees_din <= x"68fec904";
		wait for Clk_period;
		Addr <=  "0011001010111";
		Trees_din <= x"fff61995";
		wait for Clk_period;
		Addr <=  "0011001011000";
		Trees_din <= x"00691995";
		wait for Clk_period;
		Addr <=  "0011001011001";
		Trees_din <= x"9cff0e08";
		wait for Clk_period;
		Addr <=  "0011001011010";
		Trees_din <= x"da004f04";
		wait for Clk_period;
		Addr <=  "0011001011011";
		Trees_din <= x"fffd1995";
		wait for Clk_period;
		Addr <=  "0011001011100";
		Trees_din <= x"00531995";
		wait for Clk_period;
		Addr <=  "0011001011101";
		Trees_din <= x"a3fee804";
		wait for Clk_period;
		Addr <=  "0011001011110";
		Trees_din <= x"fffe1995";
		wait for Clk_period;
		Addr <=  "0011001011111";
		Trees_din <= x"ff8a1995";
		wait for Clk_period;
		Addr <=  "0011001100000";
		Trees_din <= x"9bffe608";
		wait for Clk_period;
		Addr <=  "0011001100001";
		Trees_din <= x"0fffea04";
		wait for Clk_period;
		Addr <=  "0011001100010";
		Trees_din <= x"ff821995";
		wait for Clk_period;
		Addr <=  "0011001100011";
		Trees_din <= x"fff51995";
		wait for Clk_period;
		Addr <=  "0011001100100";
		Trees_din <= x"00361995";
		wait for Clk_period;
		Addr <=  "0011001100101";
		Trees_din <= x"9eff7834";
		wait for Clk_period;
		Addr <=  "0011001100110";
		Trees_din <= x"6bff132c";
		wait for Clk_period;
		Addr <=  "0011001100111";
		Trees_din <= x"98ff3318";
		wait for Clk_period;
		Addr <=  "0011001101000";
		Trees_din <= x"80ff7a0c";
		wait for Clk_period;
		Addr <=  "0011001101001";
		Trees_din <= x"2bfeec04";
		wait for Clk_period;
		Addr <=  "0011001101010";
		Trees_din <= x"00491a31";
		wait for Clk_period;
		Addr <=  "0011001101011";
		Trees_din <= x"f5ff7104";
		wait for Clk_period;
		Addr <=  "0011001101100";
		Trees_din <= x"fffb1a31";
		wait for Clk_period;
		Addr <=  "0011001101101";
		Trees_din <= x"ff831a31";
		wait for Clk_period;
		Addr <=  "0011001101110";
		Trees_din <= x"5bff9708";
		wait for Clk_period;
		Addr <=  "0011001101111";
		Trees_din <= x"baff8004";
		wait for Clk_period;
		Addr <=  "0011001110000";
		Trees_din <= x"ffc81a31";
		wait for Clk_period;
		Addr <=  "0011001110001";
		Trees_din <= x"00471a31";
		wait for Clk_period;
		Addr <=  "0011001110010";
		Trees_din <= x"ffb31a31";
		wait for Clk_period;
		Addr <=  "0011001110011";
		Trees_din <= x"58feaf08";
		wait for Clk_period;
		Addr <=  "0011001110100";
		Trees_din <= x"71fe8604";
		wait for Clk_period;
		Addr <=  "0011001110101";
		Trees_din <= x"002d1a31";
		wait for Clk_period;
		Addr <=  "0011001110110";
		Trees_din <= x"ffa61a31";
		wait for Clk_period;
		Addr <=  "0011001110111";
		Trees_din <= x"50ffa708";
		wait for Clk_period;
		Addr <=  "0011001111000";
		Trees_din <= x"efff1d04";
		wait for Clk_period;
		Addr <=  "0011001111001";
		Trees_din <= x"00031a31";
		wait for Clk_period;
		Addr <=  "0011001111010";
		Trees_din <= x"007b1a31";
		wait for Clk_period;
		Addr <=  "0011001111011";
		Trees_din <= x"ffe51a31";
		wait for Clk_period;
		Addr <=  "0011001111100";
		Trees_din <= x"3effb404";
		wait for Clk_period;
		Addr <=  "0011001111101";
		Trees_din <= x"ff8a1a31";
		wait for Clk_period;
		Addr <=  "0011001111110";
		Trees_din <= x"00131a31";
		wait for Clk_period;
		Addr <=  "0011001111111";
		Trees_din <= x"23ff9e18";
		wait for Clk_period;
		Addr <=  "0011010000000";
		Trees_din <= x"baff6208";
		wait for Clk_period;
		Addr <=  "0011010000001";
		Trees_din <= x"0cfe8404";
		wait for Clk_period;
		Addr <=  "0011010000010";
		Trees_din <= x"006b1a31";
		wait for Clk_period;
		Addr <=  "0011010000011";
		Trees_din <= x"ffbe1a31";
		wait for Clk_period;
		Addr <=  "0011010000100";
		Trees_din <= x"1cffbc08";
		wait for Clk_period;
		Addr <=  "0011010000101";
		Trees_din <= x"52fecd04";
		wait for Clk_period;
		Addr <=  "0011010000110";
		Trees_din <= x"ffff1a31";
		wait for Clk_period;
		Addr <=  "0011010000111";
		Trees_din <= x"ff811a31";
		wait for Clk_period;
		Addr <=  "0011010001000";
		Trees_din <= x"b7ff5904";
		wait for Clk_period;
		Addr <=  "0011010001001";
		Trees_din <= x"004d1a31";
		wait for Clk_period;
		Addr <=  "0011010001010";
		Trees_din <= x"ffe01a31";
		wait for Clk_period;
		Addr <=  "0011010001011";
		Trees_din <= x"ff801a31";
		wait for Clk_period;
		Addr <=  "0011010001100";
		Trees_din <= x"b4ff6f48";
		wait for Clk_period;
		Addr <=  "0011010001101";
		Trees_din <= x"58fea910";
		wait for Clk_period;
		Addr <=  "0011010001110";
		Trees_din <= x"73004508";
		wait for Clk_period;
		Addr <=  "0011010001111";
		Trees_din <= x"71fe8604";
		wait for Clk_period;
		Addr <=  "0011010010000";
		Trees_din <= x"fffd1acd";
		wait for Clk_period;
		Addr <=  "0011010010001";
		Trees_din <= x"ff7f1acd";
		wait for Clk_period;
		Addr <=  "0011010010010";
		Trees_din <= x"6bfee604";
		wait for Clk_period;
		Addr <=  "0011010010011";
		Trees_din <= x"ffe21acd";
		wait for Clk_period;
		Addr <=  "0011010010100";
		Trees_din <= x"00571acd";
		wait for Clk_period;
		Addr <=  "0011010010101";
		Trees_din <= x"79ff131c";
		wait for Clk_period;
		Addr <=  "0011010010110";
		Trees_din <= x"46fee210";
		wait for Clk_period;
		Addr <=  "0011010010111";
		Trees_din <= x"17ffd808";
		wait for Clk_period;
		Addr <=  "0011010011000";
		Trees_din <= x"9eff4a04";
		wait for Clk_period;
		Addr <=  "0011010011001";
		Trees_din <= x"00501acd";
		wait for Clk_period;
		Addr <=  "0011010011010";
		Trees_din <= x"fff91acd";
		wait for Clk_period;
		Addr <=  "0011010011011";
		Trees_din <= x"31005504";
		wait for Clk_period;
		Addr <=  "0011010011100";
		Trees_din <= x"ff9a1acd";
		wait for Clk_period;
		Addr <=  "0011010011101";
		Trees_din <= x"00231acd";
		wait for Clk_period;
		Addr <=  "0011010011110";
		Trees_din <= x"9fff9a08";
		wait for Clk_period;
		Addr <=  "0011010011111";
		Trees_din <= x"eeff9c04";
		wait for Clk_period;
		Addr <=  "0011010100000";
		Trees_din <= x"fff81acd";
		wait for Clk_period;
		Addr <=  "0011010100001";
		Trees_din <= x"00741acd";
		wait for Clk_period;
		Addr <=  "0011010100010";
		Trees_din <= x"ffec1acd";
		wait for Clk_period;
		Addr <=  "0011010100011";
		Trees_din <= x"0700250c";
		wait for Clk_period;
		Addr <=  "0011010100100";
		Trees_din <= x"deffc108";
		wait for Clk_period;
		Addr <=  "0011010100101";
		Trees_din <= x"4afed804";
		wait for Clk_period;
		Addr <=  "0011010100110";
		Trees_din <= x"00431acd";
		wait for Clk_period;
		Addr <=  "0011010100111";
		Trees_din <= x"ffc21acd";
		wait for Clk_period;
		Addr <=  "0011010101000";
		Trees_din <= x"ff831acd";
		wait for Clk_period;
		Addr <=  "0011010101001";
		Trees_din <= x"db000908";
		wait for Clk_period;
		Addr <=  "0011010101010";
		Trees_din <= x"44000604";
		wait for Clk_period;
		Addr <=  "0011010101011";
		Trees_din <= x"ffea1acd";
		wait for Clk_period;
		Addr <=  "0011010101100";
		Trees_din <= x"005f1acd";
		wait for Clk_period;
		Addr <=  "0011010101101";
		Trees_din <= x"15ffe304";
		wait for Clk_period;
		Addr <=  "0011010101110";
		Trees_din <= x"ffab1acd";
		wait for Clk_period;
		Addr <=  "0011010101111";
		Trees_din <= x"00151acd";
		wait for Clk_period;
		Addr <=  "0011010110000";
		Trees_din <= x"d1ff8b04";
		wait for Clk_period;
		Addr <=  "0011010110001";
		Trees_din <= x"ff8a1acd";
		wait for Clk_period;
		Addr <=  "0011010110010";
		Trees_din <= x"fffe1acd";
		wait for Clk_period;
		Addr <=  "0011010110011";
		Trees_din <= x"42ff892c";
		wait for Clk_period;
		Addr <=  "0011010110100";
		Trees_din <= x"44ffb90c";
		wait for Clk_period;
		Addr <=  "0011010110101";
		Trees_din <= x"8a004308";
		wait for Clk_period;
		Addr <=  "0011010110110";
		Trees_din <= x"10003d04";
		wait for Clk_period;
		Addr <=  "0011010110111";
		Trees_din <= x"ff861b59";
		wait for Clk_period;
		Addr <=  "0011010111000";
		Trees_din <= x"ffef1b59";
		wait for Clk_period;
		Addr <=  "0011010111001";
		Trees_din <= x"00271b59";
		wait for Clk_period;
		Addr <=  "0011010111010";
		Trees_din <= x"0bff8808";
		wait for Clk_period;
		Addr <=  "0011010111011";
		Trees_din <= x"4bfe1d04";
		wait for Clk_period;
		Addr <=  "0011010111100";
		Trees_din <= x"00301b59";
		wait for Clk_period;
		Addr <=  "0011010111101";
		Trees_din <= x"ff9c1b59";
		wait for Clk_period;
		Addr <=  "0011010111110";
		Trees_din <= x"58fea908";
		wait for Clk_period;
		Addr <=  "0011010111111";
		Trees_din <= x"d4fee004";
		wait for Clk_period;
		Addr <=  "0011011000000";
		Trees_din <= x"00301b59";
		wait for Clk_period;
		Addr <=  "0011011000001";
		Trees_din <= x"ff981b59";
		wait for Clk_period;
		Addr <=  "0011011000010";
		Trees_din <= x"46fecc08";
		wait for Clk_period;
		Addr <=  "0011011000011";
		Trees_din <= x"17ffe504";
		wait for Clk_period;
		Addr <=  "0011011000100";
		Trees_din <= x"00331b59";
		wait for Clk_period;
		Addr <=  "0011011000101";
		Trees_din <= x"ffa01b59";
		wait for Clk_period;
		Addr <=  "0011011000110";
		Trees_din <= x"c8ffb304";
		wait for Clk_period;
		Addr <=  "0011011000111";
		Trees_din <= x"ffe21b59";
		wait for Clk_period;
		Addr <=  "0011011001000";
		Trees_din <= x"00521b59";
		wait for Clk_period;
		Addr <=  "0011011001001";
		Trees_din <= x"4afe9608";
		wait for Clk_period;
		Addr <=  "0011011001010";
		Trees_din <= x"1f001504";
		wait for Clk_period;
		Addr <=  "0011011001011";
		Trees_din <= x"ffe61b59";
		wait for Clk_period;
		Addr <=  "0011011001100";
		Trees_din <= x"00531b59";
		wait for Clk_period;
		Addr <=  "0011011001101";
		Trees_din <= x"92fe8f08";
		wait for Clk_period;
		Addr <=  "0011011001110";
		Trees_din <= x"c1fee904";
		wait for Clk_period;
		Addr <=  "0011011001111";
		Trees_din <= x"ffc81b59";
		wait for Clk_period;
		Addr <=  "0011011010000";
		Trees_din <= x"00481b59";
		wait for Clk_period;
		Addr <=  "0011011010001";
		Trees_din <= x"b1fe9204";
		wait for Clk_period;
		Addr <=  "0011011010010";
		Trees_din <= x"000c1b59";
		wait for Clk_period;
		Addr <=  "0011011010011";
		Trees_din <= x"1f00a904";
		wait for Clk_period;
		Addr <=  "0011011010100";
		Trees_din <= x"ff781b59";
		wait for Clk_period;
		Addr <=  "0011011010101";
		Trees_din <= x"ffe51b59";
		wait for Clk_period;
		Addr <=  "0011011010110";
		Trees_din <= x"cdff9c24";
		wait for Clk_period;
		Addr <=  "0011011010111";
		Trees_din <= x"7affe51c";
		wait for Clk_period;
		Addr <=  "0011011011000";
		Trees_din <= x"29ffa814";
		wait for Clk_period;
		Addr <=  "0011011011001";
		Trees_din <= x"baffeb0c";
		wait for Clk_period;
		Addr <=  "0011011011010";
		Trees_din <= x"5cffda04";
		wait for Clk_period;
		Addr <=  "0011011011011";
		Trees_din <= x"ffe81c0d";
		wait for Clk_period;
		Addr <=  "0011011011100";
		Trees_din <= x"7cfff704";
		wait for Clk_period;
		Addr <=  "0011011011101";
		Trees_din <= x"00711c0d";
		wait for Clk_period;
		Addr <=  "0011011011110";
		Trees_din <= x"00081c0d";
		wait for Clk_period;
		Addr <=  "0011011011111";
		Trees_din <= x"d9fffc04";
		wait for Clk_period;
		Addr <=  "0011011100000";
		Trees_din <= x"ffb91c0d";
		wait for Clk_period;
		Addr <=  "0011011100001";
		Trees_din <= x"003d1c0d";
		wait for Clk_period;
		Addr <=  "0011011100010";
		Trees_din <= x"83ff6204";
		wait for Clk_period;
		Addr <=  "0011011100011";
		Trees_din <= x"ffac1c0d";
		wait for Clk_period;
		Addr <=  "0011011100100";
		Trees_din <= x"fffe1c0d";
		wait for Clk_period;
		Addr <=  "0011011100101";
		Trees_din <= x"12003604";
		wait for Clk_period;
		Addr <=  "0011011100110";
		Trees_din <= x"ff9a1c0d";
		wait for Clk_period;
		Addr <=  "0011011100111";
		Trees_din <= x"00131c0d";
		wait for Clk_period;
		Addr <=  "0011011101000";
		Trees_din <= x"b7ff4914";
		wait for Clk_period;
		Addr <=  "0011011101001";
		Trees_din <= x"3bff5408";
		wait for Clk_period;
		Addr <=  "0011011101010";
		Trees_din <= x"2dfe7104";
		wait for Clk_period;
		Addr <=  "0011011101011";
		Trees_din <= x"002d1c0d";
		wait for Clk_period;
		Addr <=  "0011011101100";
		Trees_din <= x"ffaf1c0d";
		wait for Clk_period;
		Addr <=  "0011011101101";
		Trees_din <= x"0cfe8104";
		wait for Clk_period;
		Addr <=  "0011011101110";
		Trees_din <= x"fffc1c0d";
		wait for Clk_period;
		Addr <=  "0011011101111";
		Trees_din <= x"7affb204";
		wait for Clk_period;
		Addr <=  "0011011110000";
		Trees_din <= x"001f1c0d";
		wait for Clk_period;
		Addr <=  "0011011110001";
		Trees_din <= x"00681c0d";
		wait for Clk_period;
		Addr <=  "0011011110010";
		Trees_din <= x"d0004814";
		wait for Clk_period;
		Addr <=  "0011011110011";
		Trees_din <= x"3cfef00c";
		wait for Clk_period;
		Addr <=  "0011011110100";
		Trees_din <= x"e7ff6708";
		wait for Clk_period;
		Addr <=  "0011011110101";
		Trees_din <= x"5a00d704";
		wait for Clk_period;
		Addr <=  "0011011110110";
		Trees_din <= x"00151c0d";
		wait for Clk_period;
		Addr <=  "0011011110111";
		Trees_din <= x"00701c0d";
		wait for Clk_period;
		Addr <=  "0011011111000";
		Trees_din <= x"ffde1c0d";
		wait for Clk_period;
		Addr <=  "0011011111001";
		Trees_din <= x"00fef104";
		wait for Clk_period;
		Addr <=  "0011011111010";
		Trees_din <= x"00251c0d";
		wait for Clk_period;
		Addr <=  "0011011111011";
		Trees_din <= x"ff911c0d";
		wait for Clk_period;
		Addr <=  "0011011111100";
		Trees_din <= x"9efef704";
		wait for Clk_period;
		Addr <=  "0011011111101";
		Trees_din <= x"00181c0d";
		wait for Clk_period;
		Addr <=  "0011011111110";
		Trees_din <= x"f0fea304";
		wait for Clk_period;
		Addr <=  "0011011111111";
		Trees_din <= x"fffc1c0d";
		wait for Clk_period;
		Addr <=  "0011100000000";
		Trees_din <= x"5affef04";
		wait for Clk_period;
		Addr <=  "0011100000001";
		Trees_din <= x"ffdd1c0d";
		wait for Clk_period;
		Addr <=  "0011100000010";
		Trees_din <= x"ff761c0d";
		wait for Clk_period;
		Addr <=  "0011100000011";
		Trees_din <= x"25ffd70c";
		wait for Clk_period;
		Addr <=  "0011100000100";
		Trees_din <= x"e7ff2308";
		wait for Clk_period;
		Addr <=  "0011100000101";
		Trees_din <= x"43ffbf04";
		wait for Clk_period;
		Addr <=  "0011100000110";
		Trees_din <= x"ffd31ca1";
		wait for Clk_period;
		Addr <=  "0011100000111";
		Trees_din <= x"00461ca1";
		wait for Clk_period;
		Addr <=  "0011100001000";
		Trees_din <= x"ff8c1ca1";
		wait for Clk_period;
		Addr <=  "0011100001001";
		Trees_din <= x"98ff3328";
		wait for Clk_period;
		Addr <=  "0011100001010";
		Trees_din <= x"44002f14";
		wait for Clk_period;
		Addr <=  "0011100001011";
		Trees_din <= x"62ff2910";
		wait for Clk_period;
		Addr <=  "0011100001100";
		Trees_din <= x"f5ffac08";
		wait for Clk_period;
		Addr <=  "0011100001101";
		Trees_din <= x"c3fff204";
		wait for Clk_period;
		Addr <=  "0011100001110";
		Trees_din <= x"004d1ca1";
		wait for Clk_period;
		Addr <=  "0011100001111";
		Trees_din <= x"fff01ca1";
		wait for Clk_period;
		Addr <=  "0011100010000";
		Trees_din <= x"68ff2a04";
		wait for Clk_period;
		Addr <=  "0011100010001";
		Trees_din <= x"ff9c1ca1";
		wait for Clk_period;
		Addr <=  "0011100010010";
		Trees_din <= x"000a1ca1";
		wait for Clk_period;
		Addr <=  "0011100010011";
		Trees_din <= x"ff871ca1";
		wait for Clk_period;
		Addr <=  "0011100010100";
		Trees_din <= x"8dfe920c";
		wait for Clk_period;
		Addr <=  "0011100010101";
		Trees_din <= x"24ff5f04";
		wait for Clk_period;
		Addr <=  "0011100010110";
		Trees_din <= x"ffc81ca1";
		wait for Clk_period;
		Addr <=  "0011100010111";
		Trees_din <= x"9cff5c04";
		wait for Clk_period;
		Addr <=  "0011100011000";
		Trees_din <= x"006f1ca1";
		wait for Clk_period;
		Addr <=  "0011100011001";
		Trees_din <= x"fffc1ca1";
		wait for Clk_period;
		Addr <=  "0011100011010";
		Trees_din <= x"e6ffff04";
		wait for Clk_period;
		Addr <=  "0011100011011";
		Trees_din <= x"ffa91ca1";
		wait for Clk_period;
		Addr <=  "0011100011100";
		Trees_din <= x"002e1ca1";
		wait for Clk_period;
		Addr <=  "0011100011101";
		Trees_din <= x"a2ffcc10";
		wait for Clk_period;
		Addr <=  "0011100011110";
		Trees_din <= x"0affd504";
		wait for Clk_period;
		Addr <=  "0011100011111";
		Trees_din <= x"ffde1ca1";
		wait for Clk_period;
		Addr <=  "0011100100000";
		Trees_din <= x"2dff1608";
		wait for Clk_period;
		Addr <=  "0011100100001";
		Trees_din <= x"29ff9704";
		wait for Clk_period;
		Addr <=  "0011100100010";
		Trees_din <= x"00721ca1";
		wait for Clk_period;
		Addr <=  "0011100100011";
		Trees_din <= x"000a1ca1";
		wait for Clk_period;
		Addr <=  "0011100100100";
		Trees_din <= x"fff41ca1";
		wait for Clk_period;
		Addr <=  "0011100100101";
		Trees_din <= x"5fff5204";
		wait for Clk_period;
		Addr <=  "0011100100110";
		Trees_din <= x"ffb11ca1";
		wait for Clk_period;
		Addr <=  "0011100100111";
		Trees_din <= x"00081ca1";
		wait for Clk_period;
		Addr <=  "0011100101000";
		Trees_din <= x"15ffaa28";
		wait for Clk_period;
		Addr <=  "0011100101001";
		Trees_din <= x"fbff1308";
		wait for Clk_period;
		Addr <=  "0011100101010";
		Trees_din <= x"87ff9104";
		wait for Clk_period;
		Addr <=  "0011100101011";
		Trees_din <= x"fff71d35";
		wait for Clk_period;
		Addr <=  "0011100101100";
		Trees_din <= x"005d1d35";
		wait for Clk_period;
		Addr <=  "0011100101101";
		Trees_din <= x"da005514";
		wait for Clk_period;
		Addr <=  "0011100101110";
		Trees_din <= x"bffec208";
		wait for Clk_period;
		Addr <=  "0011100101111";
		Trees_din <= x"2fff0404";
		wait for Clk_period;
		Addr <=  "0011100110000";
		Trees_din <= x"00381d35";
		wait for Clk_period;
		Addr <=  "0011100110001";
		Trees_din <= x"ffd31d35";
		wait for Clk_period;
		Addr <=  "0011100110010";
		Trees_din <= x"5c00ea08";
		wait for Clk_period;
		Addr <=  "0011100110011";
		Trees_din <= x"dc008c04";
		wait for Clk_period;
		Addr <=  "0011100110100";
		Trees_din <= x"ff7f1d35";
		wait for Clk_period;
		Addr <=  "0011100110101";
		Trees_din <= x"fff71d35";
		wait for Clk_period;
		Addr <=  "0011100110110";
		Trees_din <= x"001d1d35";
		wait for Clk_period;
		Addr <=  "0011100110111";
		Trees_din <= x"82ff6f04";
		wait for Clk_period;
		Addr <=  "0011100111000";
		Trees_din <= x"ffc81d35";
		wait for Clk_period;
		Addr <=  "0011100111001";
		Trees_din <= x"cb002a04";
		wait for Clk_period;
		Addr <=  "0011100111010";
		Trees_din <= x"ffff1d35";
		wait for Clk_period;
		Addr <=  "0011100111011";
		Trees_din <= x"00601d35";
		wait for Clk_period;
		Addr <=  "0011100111100";
		Trees_din <= x"03ff3d08";
		wait for Clk_period;
		Addr <=  "0011100111101";
		Trees_din <= x"37ffd904";
		wait for Clk_period;
		Addr <=  "0011100111110";
		Trees_din <= x"ffa21d35";
		wait for Clk_period;
		Addr <=  "0011100111111";
		Trees_din <= x"00041d35";
		wait for Clk_period;
		Addr <=  "0011101000000";
		Trees_din <= x"87ff8c14";
		wait for Clk_period;
		Addr <=  "0011101000001";
		Trees_din <= x"46fec908";
		wait for Clk_period;
		Addr <=  "0011101000010";
		Trees_din <= x"6d005f04";
		wait for Clk_period;
		Addr <=  "0011101000011";
		Trees_din <= x"ffa61d35";
		wait for Clk_period;
		Addr <=  "0011101000100";
		Trees_din <= x"002f1d35";
		wait for Clk_period;
		Addr <=  "0011101000101";
		Trees_din <= x"c0ff9908";
		wait for Clk_period;
		Addr <=  "0011101000110";
		Trees_din <= x"7afff804";
		wait for Clk_period;
		Addr <=  "0011101000111";
		Trees_din <= x"00571d35";
		wait for Clk_period;
		Addr <=  "0011101001000";
		Trees_din <= x"ffe71d35";
		wait for Clk_period;
		Addr <=  "0011101001001";
		Trees_din <= x"ffde1d35";
		wait for Clk_period;
		Addr <=  "0011101001010";
		Trees_din <= x"6a000404";
		wait for Clk_period;
		Addr <=  "0011101001011";
		Trees_din <= x"ff9f1d35";
		wait for Clk_period;
		Addr <=  "0011101001100";
		Trees_din <= x"003c1d35";
		wait for Clk_period;
		Addr <=  "0011101001101";
		Trees_din <= x"79ff1320";
		wait for Clk_period;
		Addr <=  "0011101001110";
		Trees_din <= x"1300be0c";
		wait for Clk_period;
		Addr <=  "0011101001111";
		Trees_din <= x"c7fea308";
		wait for Clk_period;
		Addr <=  "0011101010000";
		Trees_din <= x"d7005904";
		wait for Clk_period;
		Addr <=  "0011101010001";
		Trees_din <= x"003c1dd1";
		wait for Clk_period;
		Addr <=  "0011101010010";
		Trees_din <= x"ffdc1dd1";
		wait for Clk_period;
		Addr <=  "0011101010011";
		Trees_din <= x"ffa31dd1";
		wait for Clk_period;
		Addr <=  "0011101010100";
		Trees_din <= x"50ffa310";
		wait for Clk_period;
		Addr <=  "0011101010101";
		Trees_din <= x"7dff8204";
		wait for Clk_period;
		Addr <=  "0011101010110";
		Trees_din <= x"ffe31dd1";
		wait for Clk_period;
		Addr <=  "0011101010111";
		Trees_din <= x"eeff9e04";
		wait for Clk_period;
		Addr <=  "0011101011000";
		Trees_din <= x"fffc1dd1";
		wait for Clk_period;
		Addr <=  "0011101011001";
		Trees_din <= x"b4fef904";
		wait for Clk_period;
		Addr <=  "0011101011010";
		Trees_din <= x"00731dd1";
		wait for Clk_period;
		Addr <=  "0011101011011";
		Trees_din <= x"00161dd1";
		wait for Clk_period;
		Addr <=  "0011101011100";
		Trees_din <= x"ffc91dd1";
		wait for Clk_period;
		Addr <=  "0011101011101";
		Trees_din <= x"adff661c";
		wait for Clk_period;
		Addr <=  "0011101011110";
		Trees_din <= x"b7ff7910";
		wait for Clk_period;
		Addr <=  "0011101011111";
		Trees_din <= x"58ff2c08";
		wait for Clk_period;
		Addr <=  "0011101100000";
		Trees_din <= x"65ffb904";
		wait for Clk_period;
		Addr <=  "0011101100001";
		Trees_din <= x"ffc51dd1";
		wait for Clk_period;
		Addr <=  "0011101100010";
		Trees_din <= x"002e1dd1";
		wait for Clk_period;
		Addr <=  "0011101100011";
		Trees_din <= x"29ff3604";
		wait for Clk_period;
		Addr <=  "0011101100100";
		Trees_din <= x"006a1dd1";
		wait for Clk_period;
		Addr <=  "0011101100101";
		Trees_din <= x"00021dd1";
		wait for Clk_period;
		Addr <=  "0011101100110";
		Trees_din <= x"12007008";
		wait for Clk_period;
		Addr <=  "0011101100111";
		Trees_din <= x"22ffe304";
		wait for Clk_period;
		Addr <=  "0011101101000";
		Trees_din <= x"00091dd1";
		wait for Clk_period;
		Addr <=  "0011101101001";
		Trees_din <= x"ff921dd1";
		wait for Clk_period;
		Addr <=  "0011101101010";
		Trees_din <= x"00311dd1";
		wait for Clk_period;
		Addr <=  "0011101101011";
		Trees_din <= x"f6ff4c0c";
		wait for Clk_period;
		Addr <=  "0011101101100";
		Trees_din <= x"15001508";
		wait for Clk_period;
		Addr <=  "0011101101101";
		Trees_din <= x"edff5304";
		wait for Clk_period;
		Addr <=  "0011101101110";
		Trees_din <= x"ffe11dd1";
		wait for Clk_period;
		Addr <=  "0011101101111";
		Trees_din <= x"ff7e1dd1";
		wait for Clk_period;
		Addr <=  "0011101110000";
		Trees_din <= x"fff61dd1";
		wait for Clk_period;
		Addr <=  "0011101110001";
		Trees_din <= x"03ff6604";
		wait for Clk_period;
		Addr <=  "0011101110010";
		Trees_din <= x"004d1dd1";
		wait for Clk_period;
		Addr <=  "0011101110011";
		Trees_din <= x"ffc11dd1";
		wait for Clk_period;
		Addr <=  "0011101110100";
		Trees_din <= x"25001918";
		wait for Clk_period;
		Addr <=  "0011101110101";
		Trees_din <= x"28feaf08";
		wait for Clk_period;
		Addr <=  "0011101110110";
		Trees_din <= x"35fe9204";
		wait for Clk_period;
		Addr <=  "0011101110111";
		Trees_din <= x"004c1e5d";
		wait for Clk_period;
		Addr <=  "0011101111000";
		Trees_din <= x"ffe01e5d";
		wait for Clk_period;
		Addr <=  "0011101111001";
		Trees_din <= x"68fe2f04";
		wait for Clk_period;
		Addr <=  "0011101111010";
		Trees_din <= x"00311e5d";
		wait for Clk_period;
		Addr <=  "0011101111011";
		Trees_din <= x"0b005208";
		wait for Clk_period;
		Addr <=  "0011101111100";
		Trees_din <= x"1dff7704";
		wait for Clk_period;
		Addr <=  "0011101111101";
		Trees_din <= x"ff7f1e5d";
		wait for Clk_period;
		Addr <=  "0011101111110";
		Trees_din <= x"ffdb1e5d";
		wait for Clk_period;
		Addr <=  "0011101111111";
		Trees_din <= x"00021e5d";
		wait for Clk_period;
		Addr <=  "0011110000000";
		Trees_din <= x"4aff4928";
		wait for Clk_period;
		Addr <=  "0011110000001";
		Trees_din <= x"d1ff4518";
		wait for Clk_period;
		Addr <=  "0011110000010";
		Trees_din <= x"9dff1b08";
		wait for Clk_period;
		Addr <=  "0011110000011";
		Trees_din <= x"49ffeb04";
		wait for Clk_period;
		Addr <=  "0011110000100";
		Trees_din <= x"005c1e5d";
		wait for Clk_period;
		Addr <=  "0011110000101";
		Trees_din <= x"00101e5d";
		wait for Clk_period;
		Addr <=  "0011110000110";
		Trees_din <= x"5dffa308";
		wait for Clk_period;
		Addr <=  "0011110000111";
		Trees_din <= x"a8ff7904";
		wait for Clk_period;
		Addr <=  "0011110001000";
		Trees_din <= x"ffb11e5d";
		wait for Clk_period;
		Addr <=  "0011110001001";
		Trees_din <= x"00341e5d";
		wait for Clk_period;
		Addr <=  "0011110001010";
		Trees_din <= x"83fed904";
		wait for Clk_period;
		Addr <=  "0011110001011";
		Trees_din <= x"ffe31e5d";
		wait for Clk_period;
		Addr <=  "0011110001100";
		Trees_din <= x"ff911e5d";
		wait for Clk_period;
		Addr <=  "0011110001101";
		Trees_din <= x"b7ffbf0c";
		wait for Clk_period;
		Addr <=  "0011110001110";
		Trees_din <= x"a7ffee08";
		wait for Clk_period;
		Addr <=  "0011110001111";
		Trees_din <= x"87ff6d04";
		wait for Clk_period;
		Addr <=  "0011110010000";
		Trees_din <= x"006d1e5d";
		wait for Clk_period;
		Addr <=  "0011110010001";
		Trees_din <= x"00171e5d";
		wait for Clk_period;
		Addr <=  "0011110010010";
		Trees_din <= x"ffe81e5d";
		wait for Clk_period;
		Addr <=  "0011110010011";
		Trees_din <= x"ffca1e5d";
		wait for Clk_period;
		Addr <=  "0011110010100";
		Trees_din <= x"5dffef04";
		wait for Clk_period;
		Addr <=  "0011110010101";
		Trees_din <= x"ff981e5d";
		wait for Clk_period;
		Addr <=  "0011110010110";
		Trees_din <= x"000f1e5d";
		wait for Clk_period;
		Addr <=  "0011110010111";
		Trees_din <= x"9eff7820";
		wait for Clk_period;
		Addr <=  "0011110011000";
		Trees_din <= x"6bff1318";
		wait for Clk_period;
		Addr <=  "0011110011001";
		Trees_din <= x"c0ffa814";
		wait for Clk_period;
		Addr <=  "0011110011010";
		Trees_din <= x"c0ff1908";
		wait for Clk_period;
		Addr <=  "0011110011011";
		Trees_din <= x"15ffd704";
		wait for Clk_period;
		Addr <=  "0011110011100";
		Trees_din <= x"ffb11ec9";
		wait for Clk_period;
		Addr <=  "0011110011101";
		Trees_din <= x"00161ec9";
		wait for Clk_period;
		Addr <=  "0011110011110";
		Trees_din <= x"3effa708";
		wait for Clk_period;
		Addr <=  "0011110011111";
		Trees_din <= x"9bfebf04";
		wait for Clk_period;
		Addr <=  "0011110100000";
		Trees_din <= x"ffd61ec9";
		wait for Clk_period;
		Addr <=  "0011110100001";
		Trees_din <= x"00411ec9";
		wait for Clk_period;
		Addr <=  "0011110100010";
		Trees_din <= x"ffd31ec9";
		wait for Clk_period;
		Addr <=  "0011110100011";
		Trees_din <= x"ffc01ec9";
		wait for Clk_period;
		Addr <=  "0011110100100";
		Trees_din <= x"31ff7d04";
		wait for Clk_period;
		Addr <=  "0011110100101";
		Trees_din <= x"fff31ec9";
		wait for Clk_period;
		Addr <=  "0011110100110";
		Trees_din <= x"ffaa1ec9";
		wait for Clk_period;
		Addr <=  "0011110100111";
		Trees_din <= x"23ff9e14";
		wait for Clk_period;
		Addr <=  "0011110101000";
		Trees_din <= x"46fef104";
		wait for Clk_period;
		Addr <=  "0011110101001";
		Trees_din <= x"ffb71ec9";
		wait for Clk_period;
		Addr <=  "0011110101010";
		Trees_din <= x"52ff690c";
		wait for Clk_period;
		Addr <=  "0011110101011";
		Trees_din <= x"d3fef604";
		wait for Clk_period;
		Addr <=  "0011110101100";
		Trees_din <= x"ffea1ec9";
		wait for Clk_period;
		Addr <=  "0011110101101";
		Trees_din <= x"f4fefa04";
		wait for Clk_period;
		Addr <=  "0011110101110";
		Trees_din <= x"00111ec9";
		wait for Clk_period;
		Addr <=  "0011110101111";
		Trees_din <= x"005f1ec9";
		wait for Clk_period;
		Addr <=  "0011110110000";
		Trees_din <= x"ffc21ec9";
		wait for Clk_period;
		Addr <=  "0011110110001";
		Trees_din <= x"ff901ec9";
		wait for Clk_period;
		Addr <=  "0011110110010";
		Trees_din <= x"29ff7928";
		wait for Clk_period;
		Addr <=  "0011110110011";
		Trees_din <= x"58fed00c";
		wait for Clk_period;
		Addr <=  "0011110110100";
		Trees_din <= x"7fff7e04";
		wait for Clk_period;
		Addr <=  "0011110110101";
		Trees_din <= x"ffa61f45";
		wait for Clk_period;
		Addr <=  "0011110110110";
		Trees_din <= x"d000ed04";
		wait for Clk_period;
		Addr <=  "0011110110111";
		Trees_din <= x"ffd91f45";
		wait for Clk_period;
		Addr <=  "0011110111000";
		Trees_din <= x"003a1f45";
		wait for Clk_period;
		Addr <=  "0011110111001";
		Trees_din <= x"3bff1908";
		wait for Clk_period;
		Addr <=  "0011110111010";
		Trees_din <= x"deffc204";
		wait for Clk_period;
		Addr <=  "0011110111011";
		Trees_din <= x"001e1f45";
		wait for Clk_period;
		Addr <=  "0011110111100";
		Trees_din <= x"ffb41f45";
		wait for Clk_period;
		Addr <=  "0011110111101";
		Trees_din <= x"91ffd00c";
		wait for Clk_period;
		Addr <=  "0011110111110";
		Trees_din <= x"abffe004";
		wait for Clk_period;
		Addr <=  "0011110111111";
		Trees_din <= x"ffe81f45";
		wait for Clk_period;
		Addr <=  "0011111000000";
		Trees_din <= x"e3feed04";
		wait for Clk_period;
		Addr <=  "0011111000001";
		Trees_din <= x"00531f45";
		wait for Clk_period;
		Addr <=  "0011111000010";
		Trees_din <= x"ffec1f45";
		wait for Clk_period;
		Addr <=  "0011111000011";
		Trees_din <= x"78fef204";
		wait for Clk_period;
		Addr <=  "0011111000100";
		Trees_din <= x"002d1f45";
		wait for Clk_period;
		Addr <=  "0011111000101";
		Trees_din <= x"ffb81f45";
		wait for Clk_period;
		Addr <=  "0011111000110";
		Trees_din <= x"27000508";
		wait for Clk_period;
		Addr <=  "0011111000111";
		Trees_din <= x"8a001e04";
		wait for Clk_period;
		Addr <=  "0011111001000";
		Trees_din <= x"ff8a1f45";
		wait for Clk_period;
		Addr <=  "0011111001001";
		Trees_din <= x"fff41f45";
		wait for Clk_period;
		Addr <=  "0011111001010";
		Trees_din <= x"8effd104";
		wait for Clk_period;
		Addr <=  "0011111001011";
		Trees_din <= x"ffbb1f45";
		wait for Clk_period;
		Addr <=  "0011111001100";
		Trees_din <= x"46fee904";
		wait for Clk_period;
		Addr <=  "0011111001101";
		Trees_din <= x"ffd41f45";
		wait for Clk_period;
		Addr <=  "0011111001110";
		Trees_din <= x"c8000a04";
		wait for Clk_period;
		Addr <=  "0011111001111";
		Trees_din <= x"fff91f45";
		wait for Clk_period;
		Addr <=  "0011111010000";
		Trees_din <= x"00551f45";
		wait for Clk_period;
		Addr <=  "0011111010001";
		Trees_din <= x"4afeda20";
		wait for Clk_period;
		Addr <=  "0011111010010";
		Trees_din <= x"34001414";
		wait for Clk_period;
		Addr <=  "0011111010011";
		Trees_din <= x"45fee408";
		wait for Clk_period;
		Addr <=  "0011111010100";
		Trees_din <= x"8bffee04";
		wait for Clk_period;
		Addr <=  "0011111010101";
		Trees_din <= x"002d1fc1";
		wait for Clk_period;
		Addr <=  "0011111010110";
		Trees_din <= x"ffca1fc1";
		wait for Clk_period;
		Addr <=  "0011111010111";
		Trees_din <= x"06ff6b04";
		wait for Clk_period;
		Addr <=  "0011111011000";
		Trees_din <= x"00011fc1";
		wait for Clk_period;
		Addr <=  "0011111011001";
		Trees_din <= x"0afff904";
		wait for Clk_period;
		Addr <=  "0011111011010";
		Trees_din <= x"001a1fc1";
		wait for Clk_period;
		Addr <=  "0011111011011";
		Trees_din <= x"00671fc1";
		wait for Clk_period;
		Addr <=  "0011111011100";
		Trees_din <= x"ce000208";
		wait for Clk_period;
		Addr <=  "0011111011101";
		Trees_din <= x"b1fed204";
		wait for Clk_period;
		Addr <=  "0011111011110";
		Trees_din <= x"fffa1fc1";
		wait for Clk_period;
		Addr <=  "0011111011111";
		Trees_din <= x"ffa11fc1";
		wait for Clk_period;
		Addr <=  "0011111100000";
		Trees_din <= x"00281fc1";
		wait for Clk_period;
		Addr <=  "0011111100001";
		Trees_din <= x"42ff8d18";
		wait for Clk_period;
		Addr <=  "0011111100010";
		Trees_din <= x"3bff0904";
		wait for Clk_period;
		Addr <=  "0011111100011";
		Trees_din <= x"ffa61fc1";
		wait for Clk_period;
		Addr <=  "0011111100100";
		Trees_din <= x"19ff4208";
		wait for Clk_period;
		Addr <=  "0011111100101";
		Trees_din <= x"82ff8b04";
		wait for Clk_period;
		Addr <=  "0011111100110";
		Trees_din <= x"ffaa1fc1";
		wait for Clk_period;
		Addr <=  "0011111100111";
		Trees_din <= x"00191fc1";
		wait for Clk_period;
		Addr <=  "0011111101000";
		Trees_din <= x"f8002504";
		wait for Clk_period;
		Addr <=  "0011111101001";
		Trees_din <= x"ffdf1fc1";
		wait for Clk_period;
		Addr <=  "0011111101010";
		Trees_din <= x"29ff7104";
		wait for Clk_period;
		Addr <=  "0011111101011";
		Trees_din <= x"00531fc1";
		wait for Clk_period;
		Addr <=  "0011111101100";
		Trees_din <= x"fff71fc1";
		wait for Clk_period;
		Addr <=  "0011111101101";
		Trees_din <= x"31006404";
		wait for Clk_period;
		Addr <=  "0011111101110";
		Trees_din <= x"ff8f1fc1";
		wait for Clk_period;
		Addr <=  "0011111101111";
		Trees_din <= x"000a1fc1";
		wait for Clk_period;
		Addr <=  "0011111110000";
		Trees_din <= x"15ff8614";
		wait for Clk_period;
		Addr <=  "0011111110001";
		Trees_din <= x"6dffcd04";
		wait for Clk_period;
		Addr <=  "0011111110010";
		Trees_din <= x"002c201d";
		wait for Clk_period;
		Addr <=  "0011111110011";
		Trees_din <= x"99fe2d04";
		wait for Clk_period;
		Addr <=  "0011111110100";
		Trees_din <= x"0028201d";
		wait for Clk_period;
		Addr <=  "0011111110101";
		Trees_din <= x"bffebd04";
		wait for Clk_period;
		Addr <=  "0011111110110";
		Trees_din <= x"0003201d";
		wait for Clk_period;
		Addr <=  "0011111110111";
		Trees_din <= x"e5ff2804";
		wait for Clk_period;
		Addr <=  "0011111111000";
		Trees_din <= x"ff8b201d";
		wait for Clk_period;
		Addr <=  "0011111111001";
		Trees_din <= x"fff8201d";
		wait for Clk_period;
		Addr <=  "0011111111010";
		Trees_din <= x"64fecd04";
		wait for Clk_period;
		Addr <=  "0011111111011";
		Trees_din <= x"ffbe201d";
		wait for Clk_period;
		Addr <=  "0011111111100";
		Trees_din <= x"0bff8304";
		wait for Clk_period;
		Addr <=  "0011111111101";
		Trees_din <= x"ffcb201d";
		wait for Clk_period;
		Addr <=  "0011111111110";
		Trees_din <= x"b3feaf04";
		wait for Clk_period;
		Addr <=  "0011111111111";
		Trees_din <= x"ffd6201d";
		wait for Clk_period;
		Addr <=  "0100000000000";
		Trees_din <= x"e3fee508";
		wait for Clk_period;
		Addr <=  "0100000000001";
		Trees_din <= x"58fe9f04";
		wait for Clk_period;
		Addr <=  "0100000000010";
		Trees_din <= x"ffeb201d";
		wait for Clk_period;
		Addr <=  "0100000000011";
		Trees_din <= x"0046201d";
		wait for Clk_period;
		Addr <=  "0100000000100";
		Trees_din <= x"ebfec304";
		wait for Clk_period;
		Addr <=  "0100000000101";
		Trees_din <= x"0028201d";
		wait for Clk_period;
		Addr <=  "0100000000110";
		Trees_din <= x"ffbd201d";
		wait for Clk_period;
		Addr <=  "0100000000111";
		Trees_din <= x"98ff3328";
		wait for Clk_period;
		Addr <=  "0100000001000";
		Trees_din <= x"79ff1314";
		wait for Clk_period;
		Addr <=  "0100000001001";
		Trees_din <= x"a6ff9710";
		wait for Clk_period;
		Addr <=  "0100000001010";
		Trees_din <= x"f1ff9708";
		wait for Clk_period;
		Addr <=  "0100000001011";
		Trees_din <= x"40ffff04";
		wait for Clk_period;
		Addr <=  "0100000001100";
		Trees_din <= x"00062091";
		wait for Clk_period;
		Addr <=  "0100000001101";
		Trees_din <= x"00582091";
		wait for Clk_period;
		Addr <=  "0100000001110";
		Trees_din <= x"80ffa404";
		wait for Clk_period;
		Addr <=  "0100000001111";
		Trees_din <= x"ffc22091";
		wait for Clk_period;
		Addr <=  "0100000010000";
		Trees_din <= x"00182091";
		wait for Clk_period;
		Addr <=  "0100000010001";
		Trees_din <= x"ffb92091";
		wait for Clk_period;
		Addr <=  "0100000010010";
		Trees_din <= x"6afff30c";
		wait for Clk_period;
		Addr <=  "0100000010011";
		Trees_din <= x"9fffb008";
		wait for Clk_period;
		Addr <=  "0100000010100";
		Trees_din <= x"6d008404";
		wait for Clk_period;
		Addr <=  "0100000010101";
		Trees_din <= x"ff8b2091";
		wait for Clk_period;
		Addr <=  "0100000010110";
		Trees_din <= x"fff32091";
		wait for Clk_period;
		Addr <=  "0100000010111";
		Trees_din <= x"00022091";
		wait for Clk_period;
		Addr <=  "0100000011000";
		Trees_din <= x"4dfea404";
		wait for Clk_period;
		Addr <=  "0100000011001";
		Trees_din <= x"ffd12091";
		wait for Clk_period;
		Addr <=  "0100000011010";
		Trees_din <= x"003b2091";
		wait for Clk_period;
		Addr <=  "0100000011011";
		Trees_din <= x"a2ffc010";
		wait for Clk_period;
		Addr <=  "0100000011100";
		Trees_din <= x"e6ffe80c";
		wait for Clk_period;
		Addr <=  "0100000011101";
		Trees_din <= x"58feac04";
		wait for Clk_period;
		Addr <=  "0100000011110";
		Trees_din <= x"fffb2091";
		wait for Clk_period;
		Addr <=  "0100000011111";
		Trees_din <= x"2dff1204";
		wait for Clk_period;
		Addr <=  "0100000100000";
		Trees_din <= x"00612091";
		wait for Clk_period;
		Addr <=  "0100000100001";
		Trees_din <= x"00092091";
		wait for Clk_period;
		Addr <=  "0100000100010";
		Trees_din <= x"ffeb2091";
		wait for Clk_period;
		Addr <=  "0100000100011";
		Trees_din <= x"ffd42091";
		wait for Clk_period;
		Addr <=  "0100000100100";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  6
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"94010234";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"77002420";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"4bffff14";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"7cfe1008";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"48fed104";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"02e7009d";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"ff9c009d";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"4c00e208";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"f9fd7904";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"00a9009d";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"ff53009d";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"015c009d";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"4dff1608";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"17ff3b04";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"00ca009d";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"ff76009d";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"02d0009d";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"1cffb708";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"64ffc004";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"ff65009d";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"017b009d";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"06fed704";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"03c2009d";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"03ff4804";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"0037009d";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"ff96009d";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"1dffac0c";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"77ffe304";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"ff6b009d";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"43ff5804";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"02b9009d";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"0037009d";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"4400ad0c";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"e7ff9a08";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"54004304";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"048c009d";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"01bf009d";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"00df009d";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"ffa4009d";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"9400de3c";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"06fe4610";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"31ffda0c";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"a7fff204";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"ffee0161";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"84000704";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"02480161";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"00be0161";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"ff740161";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"77002e1c";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"4bffff10";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"7cfe1008";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"0eff0e04";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"001d0161";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"01670161";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"80009e04";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"ff580161";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"00d90161";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"96ff7904";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"ff780161";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"35feea04";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"01fe0161";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"ff9d0161";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"8cfeee08";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"1dff8004";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"ffa00161";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"01de0161";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"25004c04";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"ff710161";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"003b0161";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"1dff8708";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"b5ff4204";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"ff670161";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"01b50161";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"2eff6d08";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"34ffbc04";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"00c80161";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"ff850161";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"17ffee10";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"2a006d08";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"06ff6104";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"01e90161";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"00b30161";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"1fffbd04";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"00bb0161";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"ff910161";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"07009604";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"ff980161";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"00b70161";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"9400de40";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"06fe4614";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"31ffda10";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"5fff1608";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"f7ff4904";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"ffa90225";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"002c0225";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"e1ff5004";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"00290225";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"01950225";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"ff7a0225";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"77002e1c";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"4bffff10";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"7cfe1008";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"02ff1c04";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"00140225";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"01410225";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"80008104";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"ff5b0225";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"005d0225";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"96ff7904";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"ff7e0225";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"35feea04";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"01650225";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"ffa60225";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"8cfeee08";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"1dff8004";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"ffa80225";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"015c0225";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"f8006404";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"ff750225";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"003d0225";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"1dff8708";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"b5ff4204";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"ff6d0225";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"01500225";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"2a005a14";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"17ffee0c";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"80ff0b04";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"fffc0225";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"23ff9604";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"002d0225";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"015c0225";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"1300dc04";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"ff9b0225";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"00a10225";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"1cffe204";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"ff7e0225";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"00dd0225";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"9400de3c";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"06fe9918";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"d0002a10";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"f4ff1604";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"ff8b02d9";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"61ff7d08";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"e3fec804";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"014f02d9";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"001c02d9";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"ff9e02d9";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"59fe1e04";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"00fe02d9";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"ff6602d9";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"0200271c";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"2d003610";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"7cfe5508";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"e5fe3504";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"013402d9";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"ff8602d9";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"b0005304";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"ff5d02d9";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"000602d9";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"82fefb08";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"adff7604";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"006002d9";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"017c02d9";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"ffa002d9";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"17ffcc04";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"013f02d9";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"ffa402d9";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"b5fec208";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"1c004804";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"ff7102d9";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"00bd02d9";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"9affc014";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"1afedf0c";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"80ff0b04";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"fff502d9";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"a4000c04";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"011b02d9";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"000e02d9";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"51ff5304";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"007602d9";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"ff9302d9";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"ff9002d9";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"2bfea528";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"2dff5910";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"7cff160c";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"54000808";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"0b000104";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"00d10395";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"fffe0395";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"ff980395";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"ff6f0395";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"b5fe7504";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"ff960395";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"2eff6d04";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"ff9a0395";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"47009108";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"54006a04";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"00ff0395";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"00330395";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"1f000a04";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"00970395";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"ff9d0395";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"02ffbf20";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"7cfe3208";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"f4ff1304";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"ff9e0395";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"01130395";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"17fec808";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"16ff7104";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"ff9c0395";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"00d40395";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"48fe8a08";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"7aff3804";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"01150395";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"ff770395";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"31fe2804";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"003e0395";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"ff5e0395";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"97feed10";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"17ffcc0c";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"12007308";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"d5006a04";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"01560395";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"00580395";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"fff20395";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"ff960395";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"9c002a04";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"ff6d0395";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"00970395";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"2300742c";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"7700241c";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"2d002214";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"4bffff0c";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"44fed804";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"00780431";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"f9fd7904";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"00690431";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"ff610431";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"4dff1604";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"ff900431";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"00950431";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"c4feeb04";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"00c90431";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"ff9f0431";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"1cffb708";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"8cffb804";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"ff830431";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"00290431";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"a7000604";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"fff70431";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"00e00431";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"17ffe61c";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"2dff5208";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"7cfeb304";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"007f0431";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"ff790431";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"80ff2b08";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"f1ffbd04";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"ff950431";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"004c0431";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"b5fe5c04";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"ffac0431";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"1f005504";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"00e50431";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"004c0431";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"06fdf304";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"005f0431";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"ff6b0431";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"23007434";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"77002424";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"2d00221c";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"48fea30c";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"4dff5104";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"ff7d04e5";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"65ff6604";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"002b04e5";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"011604e5";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"02ffd908";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"17fe9e04";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"003804e5";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"ff6104e5";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"2efffa04";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"ff8304e5";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"00b504e5";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"c4feeb04";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"00b204e5";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"ffa504e5";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"d0002a0c";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"1cffb704";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"fff204e5";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"50ff3f04";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"00ca04e5";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"003304e5";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"ff8b04e5";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"17ffd920";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"1dffa10c";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"8ffe4b04";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"00be04e5";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"0eff4704";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"ff7604e5";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"003304e5";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"80ff6108";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"02ffe704";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"ff8d04e5";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"007904e5";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"a4ffee08";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"a1ffa104";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"00d504e5";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"003604e5";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"000604e5";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"06fdf304";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"008004e5";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"ff6d04e5";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"23004730";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"1c006224";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"2f00d81c";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"3000a010";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"63009e08";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"c1fdee04";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"003405b9";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"ff6305b9";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"80ffe304";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"ffab05b9";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"008e05b9";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"72ff9f04";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"00d605b9";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"f3fe9404";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"fff105b9";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"ff9605b9";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"53ff1004";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"00ad05b9";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"fffb05b9";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"80ffea08";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"aaff2404";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"fff105b9";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"ff9705b9";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"00c205b9";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"17ff6f20";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"97fefd18";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"47009110";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"80ff6108";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"72fff404";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"ffa605b9";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"008e05b9";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"88008c04";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"00d505b9";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"003605b9";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"30007104";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"ffa105b9";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"006805b9";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"e2fe5104";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"006505b9";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"ff8e05b9";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"7cfecc0c";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"b5fecd04";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"ffa405b9";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"6affb104";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"00bf05b9";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"000005b9";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"4c002308";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"2cfee704";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"fff205b9";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"ff6805b9";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"52ff1204";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"ffb305b9";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"009e05b9";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"23004738";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"1c004228";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"02ffd918";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"63009e10";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"3000ae08";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"a7013204";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"ff620685";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"fff70685";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"a6ffbc04";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"ff9f0685";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"00940685";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"80ffe304";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"ffae0685";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"00800685";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"54ffe10c";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"0fff5304";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"ffe40685";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"04002404";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"01080685";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"00460685";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"ff8a0685";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"06fefa08";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"79ff0004";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"00c00685";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"00280685";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"abffcc04";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"000c0685";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"ff840685";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"17ffef28";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"2dff500c";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"50feaa08";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"27ff9504";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"008c0685";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"fff20685";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"ff7a0685";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"f4ff4110";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"2effb108";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"06ff5804";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"ff860685";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"fff40685";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"4dff0204";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"ffc20685";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"009c0685";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"c5ff0c04";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"001b0685";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"97ff2d04";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"00bf0685";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"00110685";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"88ff6404";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"001f0685";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"ff700685";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"23004730";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"1c004220";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"02ffd914";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"3000ae0c";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"63009e08";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"a7013204";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"ff63074d";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"fff9074d";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"001c074d";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"38fefe04";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"008a074d";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"ffa3074d";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"e7ff1508";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"03ff1904";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"00d9074d";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"ffe3074d";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"ff8d074d";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"06fefa08";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"1fffe004";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"00b3074d";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"0021074d";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"1bff5004";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"000a074d";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"ff8a074d";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"17ff6f18";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"97fefd10";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"4700910c";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"81ffdb08";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"66009504";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"00bb074d";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"001a074d";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"fffc074d";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"fffd074d";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"e2fe5104";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"0056074d";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"ff99074d";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"7cfecc0c";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"b5fecd04";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"ffab074d";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"6affb104";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"00a5074d";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"fff8074d";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"4c002308";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"79fffe04";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"ff6d074d";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"ffe2074d";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"52ff1204";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"ffba074d";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"0085074d";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"06fee134";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"4dfef810";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"d0001f0c";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"f4ff4204";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"ffa807f9";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"58fee104";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"000f07f9";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"009a07f9";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"ff7607f9";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"47004a18";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"cafe0208";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"1cffd004";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"ffaa07f9";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"005707f9";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"baff4108";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"e7fea004";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"006507f9";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"ffc007f9";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"80ff5a04";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"002307f9";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"00b607f9";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"2bfe4808";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"da008b04";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"000e07f9";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"007b07f9";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"ff8e07f9";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"02ffbf14";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"2d00220c";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"17fe9e04";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"004507f9";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"24fe8704";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"003007f9";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"ff6407f9";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"0efeee04";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"ffd307f9";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"008707f9";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"97feed0c";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"4bff4b04";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"fff507f9";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"b9fed004";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"004107f9";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"00e007f9";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"ff8607f9";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"2300472c";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"06fee918";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"4dfef908";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"11ffdf04";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"ff7508a5";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"ffe408a5";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"8bffe00c";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"2a002908";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"6d002f04";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"00d508a5";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"003a08a5";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"fffd08a5";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"ffae08a5";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"02ffbf08";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"b5000b04";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"ff6508a5";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"ffee08a5";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"97feb908";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"7efed804";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"ffec08a5";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"00d208a5";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"ff8e08a5";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"17ffef24";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"b5feb308";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"17ff4a04";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"002308a5";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"ff8a08a5";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"f4ff060c";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"97febd08";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"70fecd04";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"ffc808a5";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"007c08a5";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"ff9708a5";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"50ff5008";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"a1ffb204";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"00a508a5";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"ffec08a5";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"83fee604";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"005d08a5";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"ffa708a5";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"71fe3c04";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"fffa08a5";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"ff7b08a5";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"2dff8b24";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"06feb914";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"e5fe260c";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"daffa804";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"ffe10931";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"4dff2904";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"00170931";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"009e0931";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"b6ffe504";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"ff8c0931";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"003e0931";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"02ffd908";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"6afeb504";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"fff00931";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"ff650931";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"d0000f04";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"00ac0931";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"ffae0931";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"2bff2618";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"1f005510";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"5400670c";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"aaffcf08";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"faffc504";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"00aa0931";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"00250931";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"000c0931";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"ffc60931";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"a7013204";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"ff900931";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"00460931";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"80002c08";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"39002104";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"ff740931";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"ffea0931";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"00780931";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"2dff8b24";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"06feb914";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"e5fe260c";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"bcff0904";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"ffeb09b5";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"40002004";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"001709b5";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"009909b5";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"b6ffe504";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"ff9109b5";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"003609b5";
		wait for Clk_period;
		Addr <=  "0001001010111";
		Trees_din <= x"02ffd908";
		wait for Clk_period;
		Addr <=  "0001001011000";
		Trees_din <= x"8cfe6e04";
		wait for Clk_period;
		Addr <=  "0001001011001";
		Trees_din <= x"ffe809b5";
		wait for Clk_period;
		Addr <=  "0001001011010";
		Trees_din <= x"ff6609b5";
		wait for Clk_period;
		Addr <=  "0001001011011";
		Trees_din <= x"d0000f04";
		wait for Clk_period;
		Addr <=  "0001001011100";
		Trees_din <= x"00a309b5";
		wait for Clk_period;
		Addr <=  "0001001011101";
		Trees_din <= x"ffb409b5";
		wait for Clk_period;
		Addr <=  "0001001011110";
		Trees_din <= x"17ffef18";
		wait for Clk_period;
		Addr <=  "0001001011111";
		Trees_din <= x"2bffa914";
		wait for Clk_period;
		Addr <=  "0001001100000";
		Trees_din <= x"1f00440c";
		wait for Clk_period;
		Addr <=  "0001001100001";
		Trees_din <= x"80ff5f04";
		wait for Clk_period;
		Addr <=  "0001001100010";
		Trees_din <= x"ffea09b5";
		wait for Clk_period;
		Addr <=  "0001001100011";
		Trees_din <= x"b5fec604";
		wait for Clk_period;
		Addr <=  "0001001100100";
		Trees_din <= x"000909b5";
		wait for Clk_period;
		Addr <=  "0001001100101";
		Trees_din <= x"009c09b5";
		wait for Clk_period;
		Addr <=  "0001001100110";
		Trees_din <= x"79feba04";
		wait for Clk_period;
		Addr <=  "0001001100111";
		Trees_din <= x"004009b5";
		wait for Clk_period;
		Addr <=  "0001001101000";
		Trees_din <= x"ff9709b5";
		wait for Clk_period;
		Addr <=  "0001001101001";
		Trees_din <= x"ff9509b5";
		wait for Clk_period;
		Addr <=  "0001001101010";
		Trees_din <= x"deff5004";
		wait for Clk_period;
		Addr <=  "0001001101011";
		Trees_din <= x"ffef09b5";
		wait for Clk_period;
		Addr <=  "0001001101100";
		Trees_din <= x"ff7d09b5";
		wait for Clk_period;
		Addr <=  "0001001101101";
		Trees_din <= x"06fee124";
		wait for Clk_period;
		Addr <=  "0001001101110";
		Trees_din <= x"d0003718";
		wait for Clk_period;
		Addr <=  "0001001101111";
		Trees_din <= x"4dfea708";
		wait for Clk_period;
		Addr <=  "0001001110000";
		Trees_din <= x"3eff7d04";
		wait for Clk_period;
		Addr <=  "0001001110001";
		Trees_din <= x"ffae0a31";
		wait for Clk_period;
		Addr <=  "0001001110010";
		Trees_din <= x"00380a31";
		wait for Clk_period;
		Addr <=  "0001001110011";
		Trees_din <= x"f4feb704";
		wait for Clk_period;
		Addr <=  "0001001110100";
		Trees_din <= x"ffe20a31";
		wait for Clk_period;
		Addr <=  "0001001110101";
		Trees_din <= x"cafe0204";
		wait for Clk_period;
		Addr <=  "0001001110110";
		Trees_din <= x"00070a31";
		wait for Clk_period;
		Addr <=  "0001001110111";
		Trees_din <= x"41ff6b04";
		wait for Clk_period;
		Addr <=  "0001001111000";
		Trees_din <= x"009d0a31";
		wait for Clk_period;
		Addr <=  "0001001111001";
		Trees_din <= x"00100a31";
		wait for Clk_period;
		Addr <=  "0001001111010";
		Trees_din <= x"94009c04";
		wait for Clk_period;
		Addr <=  "0001001111011";
		Trees_din <= x"ff790a31";
		wait for Clk_period;
		Addr <=  "0001001111100";
		Trees_din <= x"1dfff904";
		wait for Clk_period;
		Addr <=  "0001001111101";
		Trees_din <= x"ffd70a31";
		wait for Clk_period;
		Addr <=  "0001001111110";
		Trees_din <= x"006a0a31";
		wait for Clk_period;
		Addr <=  "0001001111111";
		Trees_din <= x"02ff900c";
		wait for Clk_period;
		Addr <=  "0001010000000";
		Trees_din <= x"17fe9e04";
		wait for Clk_period;
		Addr <=  "0001010000001";
		Trees_din <= x"00350a31";
		wait for Clk_period;
		Addr <=  "0001010000010";
		Trees_din <= x"2d002204";
		wait for Clk_period;
		Addr <=  "0001010000011";
		Trees_din <= x"ff670a31";
		wait for Clk_period;
		Addr <=  "0001010000100";
		Trees_din <= x"00240a31";
		wait for Clk_period;
		Addr <=  "0001010000101";
		Trees_din <= x"97feed0c";
		wait for Clk_period;
		Addr <=  "0001010000110";
		Trees_din <= x"4bff5504";
		wait for Clk_period;
		Addr <=  "0001010000111";
		Trees_din <= x"ffd70a31";
		wait for Clk_period;
		Addr <=  "0001010001000";
		Trees_din <= x"1cffe904";
		wait for Clk_period;
		Addr <=  "0001010001001";
		Trees_din <= x"002e0a31";
		wait for Clk_period;
		Addr <=  "0001010001010";
		Trees_din <= x"00cc0a31";
		wait for Clk_period;
		Addr <=  "0001010001011";
		Trees_din <= x"ff840a31";
		wait for Clk_period;
		Addr <=  "0001010001100";
		Trees_din <= x"23004720";
		wait for Clk_period;
		Addr <=  "0001010001101";
		Trees_din <= x"1c000210";
		wait for Clk_period;
		Addr <=  "0001010001110";
		Trees_din <= x"f9fd7904";
		wait for Clk_period;
		Addr <=  "0001010001111";
		Trees_din <= x"00500abd";
		wait for Clk_period;
		Addr <=  "0001010010000";
		Trees_din <= x"2f009a08";
		wait for Clk_period;
		Addr <=  "0001010010001";
		Trees_din <= x"4dff9504";
		wait for Clk_period;
		Addr <=  "0001010010010";
		Trees_din <= x"ff670abd";
		wait for Clk_period;
		Addr <=  "0001010010011";
		Trees_din <= x"ffe40abd";
		wait for Clk_period;
		Addr <=  "0001010010100";
		Trees_din <= x"001c0abd";
		wait for Clk_period;
		Addr <=  "0001010010101";
		Trees_din <= x"e5fe7a08";
		wait for Clk_period;
		Addr <=  "0001010010110";
		Trees_din <= x"14ff3f04";
		wait for Clk_period;
		Addr <=  "0001010010111";
		Trees_din <= x"00090abd";
		wait for Clk_period;
		Addr <=  "0001010011000";
		Trees_din <= x"00cb0abd";
		wait for Clk_period;
		Addr <=  "0001010011001";
		Trees_din <= x"2dffae04";
		wait for Clk_period;
		Addr <=  "0001010011010";
		Trees_din <= x"ff8a0abd";
		wait for Clk_period;
		Addr <=  "0001010011011";
		Trees_din <= x"00370abd";
		wait for Clk_period;
		Addr <=  "0001010011100";
		Trees_din <= x"17ff5610";
		wait for Clk_period;
		Addr <=  "0001010011101";
		Trees_din <= x"2a005a0c";
		wait for Clk_period;
		Addr <=  "0001010011110";
		Trees_din <= x"97fefd08";
		wait for Clk_period;
		Addr <=  "0001010011111";
		Trees_din <= x"24ffc704";
		wait for Clk_period;
		Addr <=  "0001010100000";
		Trees_din <= x"009c0abd";
		wait for Clk_period;
		Addr <=  "0001010100001";
		Trees_din <= x"00280abd";
		wait for Clk_period;
		Addr <=  "0001010100010";
		Trees_din <= x"ffff0abd";
		wait for Clk_period;
		Addr <=  "0001010100011";
		Trees_din <= x"ffee0abd";
		wait for Clk_period;
		Addr <=  "0001010100100";
		Trees_din <= x"e5fe0808";
		wait for Clk_period;
		Addr <=  "0001010100101";
		Trees_din <= x"27ffb404";
		wait for Clk_period;
		Addr <=  "0001010100110";
		Trees_din <= x"00760abd";
		wait for Clk_period;
		Addr <=  "0001010100111";
		Trees_din <= x"fff50abd";
		wait for Clk_period;
		Addr <=  "0001010101000";
		Trees_din <= x"e7feb408";
		wait for Clk_period;
		Addr <=  "0001010101001";
		Trees_din <= x"d7008804";
		wait for Clk_period;
		Addr <=  "0001010101010";
		Trees_din <= x"005e0abd";
		wait for Clk_period;
		Addr <=  "0001010101011";
		Trees_din <= x"fff30abd";
		wait for Clk_period;
		Addr <=  "0001010101100";
		Trees_din <= x"83fe7604";
		wait for Clk_period;
		Addr <=  "0001010101101";
		Trees_din <= x"ffda0abd";
		wait for Clk_period;
		Addr <=  "0001010101110";
		Trees_din <= x"ff7b0abd";
		wait for Clk_period;
		Addr <=  "0001010101111";
		Trees_din <= x"06fee128";
		wait for Clk_period;
		Addr <=  "0001010110000";
		Trees_din <= x"1cffbf10";
		wait for Clk_period;
		Addr <=  "0001010110001";
		Trees_din <= x"48fea308";
		wait for Clk_period;
		Addr <=  "0001010110010";
		Trees_din <= x"47ffe504";
		wait for Clk_period;
		Addr <=  "0001010110011";
		Trees_din <= x"00770b39";
		wait for Clk_period;
		Addr <=  "0001010110100";
		Trees_din <= x"ffc40b39";
		wait for Clk_period;
		Addr <=  "0001010110101";
		Trees_din <= x"21fea904";
		wait for Clk_period;
		Addr <=  "0001010110110";
		Trees_din <= x"00240b39";
		wait for Clk_period;
		Addr <=  "0001010110111";
		Trees_din <= x"ff820b39";
		wait for Clk_period;
		Addr <=  "0001010111000";
		Trees_din <= x"4dfebb08";
		wait for Clk_period;
		Addr <=  "0001010111001";
		Trees_din <= x"eeff7604";
		wait for Clk_period;
		Addr <=  "0001010111010";
		Trees_din <= x"00360b39";
		wait for Clk_period;
		Addr <=  "0001010111011";
		Trees_din <= x"ffa50b39";
		wait for Clk_period;
		Addr <=  "0001010111100";
		Trees_din <= x"73009f0c";
		wait for Clk_period;
		Addr <=  "0001010111101";
		Trees_din <= x"cafe0204";
		wait for Clk_period;
		Addr <=  "0001010111110";
		Trees_din <= x"001f0b39";
		wait for Clk_period;
		Addr <=  "0001010111111";
		Trees_din <= x"a7000304";
		wait for Clk_period;
		Addr <=  "0001011000000";
		Trees_din <= x"00250b39";
		wait for Clk_period;
		Addr <=  "0001011000001";
		Trees_din <= x"009d0b39";
		wait for Clk_period;
		Addr <=  "0001011000010";
		Trees_din <= x"fffe0b39";
		wait for Clk_period;
		Addr <=  "0001011000011";
		Trees_din <= x"02ff900c";
		wait for Clk_period;
		Addr <=  "0001011000100";
		Trees_din <= x"2dffae04";
		wait for Clk_period;
		Addr <=  "0001011000101";
		Trees_din <= x"ff680b39";
		wait for Clk_period;
		Addr <=  "0001011000110";
		Trees_din <= x"c8ffcc04";
		wait for Clk_period;
		Addr <=  "0001011000111";
		Trees_din <= x"00390b39";
		wait for Clk_period;
		Addr <=  "0001011001000";
		Trees_din <= x"ff9e0b39";
		wait for Clk_period;
		Addr <=  "0001011001001";
		Trees_din <= x"97feed08";
		wait for Clk_period;
		Addr <=  "0001011001010";
		Trees_din <= x"4bff5504";
		wait for Clk_period;
		Addr <=  "0001011001011";
		Trees_din <= x"ffdd0b39";
		wait for Clk_period;
		Addr <=  "0001011001100";
		Trees_din <= x"00a60b39";
		wait for Clk_period;
		Addr <=  "0001011001101";
		Trees_din <= x"ff8d0b39";
		wait for Clk_period;
		Addr <=  "0001011001110";
		Trees_din <= x"2300471c";
		wait for Clk_period;
		Addr <=  "0001011001111";
		Trees_din <= x"1c00020c";
		wait for Clk_period;
		Addr <=  "0001011010000";
		Trees_din <= x"2f009a08";
		wait for Clk_period;
		Addr <=  "0001011010001";
		Trees_din <= x"22ff1404";
		wait for Clk_period;
		Addr <=  "0001011010010";
		Trees_din <= x"000e0bb5";
		wait for Clk_period;
		Addr <=  "0001011010011";
		Trees_din <= x"ff690bb5";
		wait for Clk_period;
		Addr <=  "0001011010100";
		Trees_din <= x"00250bb5";
		wait for Clk_period;
		Addr <=  "0001011010101";
		Trees_din <= x"e5fe7a08";
		wait for Clk_period;
		Addr <=  "0001011010110";
		Trees_din <= x"25ffc604";
		wait for Clk_period;
		Addr <=  "0001011010111";
		Trees_din <= x"00b50bb5";
		wait for Clk_period;
		Addr <=  "0001011011000";
		Trees_din <= x"00110bb5";
		wait for Clk_period;
		Addr <=  "0001011011001";
		Trees_din <= x"2dff7104";
		wait for Clk_period;
		Addr <=  "0001011011010";
		Trees_din <= x"ff8c0bb5";
		wait for Clk_period;
		Addr <=  "0001011011011";
		Trees_din <= x"00260bb5";
		wait for Clk_period;
		Addr <=  "0001011011100";
		Trees_din <= x"f4ff4f10";
		wait for Clk_period;
		Addr <=  "0001011011101";
		Trees_din <= x"4dff5108";
		wait for Clk_period;
		Addr <=  "0001011011110";
		Trees_din <= x"da008b04";
		wait for Clk_period;
		Addr <=  "0001011011111";
		Trees_din <= x"ff850bb5";
		wait for Clk_period;
		Addr <=  "0001011100000";
		Trees_din <= x"ffed0bb5";
		wait for Clk_period;
		Addr <=  "0001011100001";
		Trees_din <= x"2effc704";
		wait for Clk_period;
		Addr <=  "0001011100010";
		Trees_din <= x"ffe90bb5";
		wait for Clk_period;
		Addr <=  "0001011100011";
		Trees_din <= x"00620bb5";
		wait for Clk_period;
		Addr <=  "0001011100100";
		Trees_din <= x"54006210";
		wait for Clk_period;
		Addr <=  "0001011100101";
		Trees_din <= x"c0ffe80c";
		wait for Clk_period;
		Addr <=  "0001011100110";
		Trees_din <= x"1dff9908";
		wait for Clk_period;
		Addr <=  "0001011100111";
		Trees_din <= x"8ffe3a04";
		wait for Clk_period;
		Addr <=  "0001011101000";
		Trees_din <= x"00590bb5";
		wait for Clk_period;
		Addr <=  "0001011101001";
		Trees_din <= x"ffe10bb5";
		wait for Clk_period;
		Addr <=  "0001011101010";
		Trees_din <= x"00930bb5";
		wait for Clk_period;
		Addr <=  "0001011101011";
		Trees_din <= x"fff80bb5";
		wait for Clk_period;
		Addr <=  "0001011101100";
		Trees_din <= x"ffcc0bb5";
		wait for Clk_period;
		Addr <=  "0001011101101";
		Trees_din <= x"06fee924";
		wait for Clk_period;
		Addr <=  "0001011101110";
		Trees_din <= x"d0003714";
		wait for Clk_period;
		Addr <=  "0001011101111";
		Trees_din <= x"1f004410";
		wait for Clk_period;
		Addr <=  "0001011110000";
		Trees_din <= x"aaffe00c";
		wait for Clk_period;
		Addr <=  "0001011110001";
		Trees_din <= x"66008008";
		wait for Clk_period;
		Addr <=  "0001011110010";
		Trees_din <= x"e4fede04";
		wait for Clk_period;
		Addr <=  "0001011110011";
		Trees_din <= x"008d0c29";
		wait for Clk_period;
		Addr <=  "0001011110100";
		Trees_din <= x"00110c29";
		wait for Clk_period;
		Addr <=  "0001011110101";
		Trees_din <= x"00060c29";
		wait for Clk_period;
		Addr <=  "0001011110110";
		Trees_din <= x"ffeb0c29";
		wait for Clk_period;
		Addr <=  "0001011110111";
		Trees_din <= x"ffea0c29";
		wait for Clk_period;
		Addr <=  "0001011111000";
		Trees_din <= x"94009c04";
		wait for Clk_period;
		Addr <=  "0001011111001";
		Trees_din <= x"ff850c29";
		wait for Clk_period;
		Addr <=  "0001011111010";
		Trees_din <= x"b3fef508";
		wait for Clk_period;
		Addr <=  "0001011111011";
		Trees_din <= x"59fe1e04";
		wait for Clk_period;
		Addr <=  "0001011111100";
		Trees_din <= x"00660c29";
		wait for Clk_period;
		Addr <=  "0001011111101";
		Trees_din <= x"000d0c29";
		wait for Clk_period;
		Addr <=  "0001011111110";
		Trees_din <= x"ffcb0c29";
		wait for Clk_period;
		Addr <=  "0001011111111";
		Trees_din <= x"02ff900c";
		wait for Clk_period;
		Addr <=  "0001100000000";
		Trees_din <= x"f4ffed08";
		wait for Clk_period;
		Addr <=  "0001100000001";
		Trees_din <= x"50fe7e04";
		wait for Clk_period;
		Addr <=  "0001100000010";
		Trees_din <= x"fff80c29";
		wait for Clk_period;
		Addr <=  "0001100000011";
		Trees_din <= x"ff690c29";
		wait for Clk_period;
		Addr <=  "0001100000100";
		Trees_din <= x"000f0c29";
		wait for Clk_period;
		Addr <=  "0001100000101";
		Trees_din <= x"97feed08";
		wait for Clk_period;
		Addr <=  "0001100000110";
		Trees_din <= x"4bff5504";
		wait for Clk_period;
		Addr <=  "0001100000111";
		Trees_din <= x"ffdc0c29";
		wait for Clk_period;
		Addr <=  "0001100001000";
		Trees_din <= x"00940c29";
		wait for Clk_period;
		Addr <=  "0001100001001";
		Trees_din <= x"ff960c29";
		wait for Clk_period;
		Addr <=  "0001100001010";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0001100001011";
		Trees_din <= x"2dff8b18";
		wait for Clk_period;
		Addr <=  "0001100001100";
		Trees_din <= x"50ff1414";
		wait for Clk_period;
		Addr <=  "0001100001101";
		Trees_din <= x"d000130c";
		wait for Clk_period;
		Addr <=  "0001100001110";
		Trees_din <= x"78ffe304";
		wait for Clk_period;
		Addr <=  "0001100001111";
		Trees_din <= x"ffd20c99";
		wait for Clk_period;
		Addr <=  "0001100010000";
		Trees_din <= x"fbff9b04";
		wait for Clk_period;
		Addr <=  "0001100010001";
		Trees_din <= x"000b0c99";
		wait for Clk_period;
		Addr <=  "0001100010010";
		Trees_din <= x"008e0c99";
		wait for Clk_period;
		Addr <=  "0001100010011";
		Trees_din <= x"94009c04";
		wait for Clk_period;
		Addr <=  "0001100010100";
		Trees_din <= x"ff7f0c99";
		wait for Clk_period;
		Addr <=  "0001100010101";
		Trees_din <= x"00210c99";
		wait for Clk_period;
		Addr <=  "0001100010110";
		Trees_din <= x"ff6c0c99";
		wait for Clk_period;
		Addr <=  "0001100010111";
		Trees_din <= x"17ffef1c";
		wait for Clk_period;
		Addr <=  "0001100011000";
		Trees_din <= x"f4feef08";
		wait for Clk_period;
		Addr <=  "0001100011001";
		Trees_din <= x"36ff4d04";
		wait for Clk_period;
		Addr <=  "0001100011010";
		Trees_din <= x"000c0c99";
		wait for Clk_period;
		Addr <=  "0001100011011";
		Trees_din <= x"ffa90c99";
		wait for Clk_period;
		Addr <=  "0001100011100";
		Trees_din <= x"a7fffb08";
		wait for Clk_period;
		Addr <=  "0001100011101";
		Trees_din <= x"f4ff8e04";
		wait for Clk_period;
		Addr <=  "0001100011110";
		Trees_din <= x"ffb60c99";
		wait for Clk_period;
		Addr <=  "0001100011111";
		Trees_din <= x"00400c99";
		wait for Clk_period;
		Addr <=  "0001100100000";
		Trees_din <= x"88005708";
		wait for Clk_period;
		Addr <=  "0001100100001";
		Trees_din <= x"b0ff0d04";
		wait for Clk_period;
		Addr <=  "0001100100010";
		Trees_din <= x"001b0c99";
		wait for Clk_period;
		Addr <=  "0001100100011";
		Trees_din <= x"008b0c99";
		wait for Clk_period;
		Addr <=  "0001100100100";
		Trees_din <= x"00050c99";
		wait for Clk_period;
		Addr <=  "0001100100101";
		Trees_din <= x"ffa00c99";
		wait for Clk_period;
		Addr <=  "0001100100110";
		Trees_din <= x"1cffd918";
		wait for Clk_period;
		Addr <=  "0001100100111";
		Trees_din <= x"7cfe3208";
		wait for Clk_period;
		Addr <=  "0001100101000";
		Trees_din <= x"e5fe0804";
		wait for Clk_period;
		Addr <=  "0001100101001";
		Trees_din <= x"005f0d05";
		wait for Clk_period;
		Addr <=  "0001100101010";
		Trees_din <= x"001a0d05";
		wait for Clk_period;
		Addr <=  "0001100101011";
		Trees_din <= x"7700240c";
		wait for Clk_period;
		Addr <=  "0001100101100";
		Trees_din <= x"80003308";
		wait for Clk_period;
		Addr <=  "0001100101101";
		Trees_din <= x"4c002304";
		wait for Clk_period;
		Addr <=  "0001100101110";
		Trees_din <= x"ff6a0d05";
		wait for Clk_period;
		Addr <=  "0001100101111";
		Trees_din <= x"ffd80d05";
		wait for Clk_period;
		Addr <=  "0001100110000";
		Trees_din <= x"fff70d05";
		wait for Clk_period;
		Addr <=  "0001100110001";
		Trees_din <= x"00130d05";
		wait for Clk_period;
		Addr <=  "0001100110010";
		Trees_din <= x"e5fe8210";
		wait for Clk_period;
		Addr <=  "0001100110011";
		Trees_din <= x"78ff8f04";
		wait for Clk_period;
		Addr <=  "0001100110100";
		Trees_din <= x"ffe10d05";
		wait for Clk_period;
		Addr <=  "0001100110101";
		Trees_din <= x"47006b08";
		wait for Clk_period;
		Addr <=  "0001100110110";
		Trees_din <= x"97fef204";
		wait for Clk_period;
		Addr <=  "0001100110111";
		Trees_din <= x"00980d05";
		wait for Clk_period;
		Addr <=  "0001100111000";
		Trees_din <= x"00200d05";
		wait for Clk_period;
		Addr <=  "0001100111001";
		Trees_din <= x"00010d05";
		wait for Clk_period;
		Addr <=  "0001100111010";
		Trees_din <= x"17ff3b08";
		wait for Clk_period;
		Addr <=  "0001100111011";
		Trees_din <= x"9400f404";
		wait for Clk_period;
		Addr <=  "0001100111100";
		Trees_din <= x"000d0d05";
		wait for Clk_period;
		Addr <=  "0001100111101";
		Trees_din <= x"00540d05";
		wait for Clk_period;
		Addr <=  "0001100111110";
		Trees_din <= x"db00e104";
		wait for Clk_period;
		Addr <=  "0001100111111";
		Trees_din <= x"ff870d05";
		wait for Clk_period;
		Addr <=  "0001101000000";
		Trees_din <= x"ffec0d05";
		wait for Clk_period;
		Addr <=  "0001101000001";
		Trees_din <= x"50ff1820";
		wait for Clk_period;
		Addr <=  "0001101000010";
		Trees_din <= x"1cffc910";
		wait for Clk_period;
		Addr <=  "0001101000011";
		Trees_din <= x"7cfecc08";
		wait for Clk_period;
		Addr <=  "0001101000100";
		Trees_din <= x"64ff3e04";
		wait for Clk_period;
		Addr <=  "0001101000101";
		Trees_din <= x"ffdb0d61";
		wait for Clk_period;
		Addr <=  "0001101000110";
		Trees_din <= x"005d0d61";
		wait for Clk_period;
		Addr <=  "0001101000111";
		Trees_din <= x"4c002304";
		wait for Clk_period;
		Addr <=  "0001101001000";
		Trees_din <= x"ff810d61";
		wait for Clk_period;
		Addr <=  "0001101001001";
		Trees_din <= x"00100d61";
		wait for Clk_period;
		Addr <=  "0001101001010";
		Trees_din <= x"17ffcc0c";
		wait for Clk_period;
		Addr <=  "0001101001011";
		Trees_din <= x"2eff9604";
		wait for Clk_period;
		Addr <=  "0001101001100";
		Trees_din <= x"fff80d61";
		wait for Clk_period;
		Addr <=  "0001101001101";
		Trees_din <= x"22fea604";
		wait for Clk_period;
		Addr <=  "0001101001110";
		Trees_din <= x"00120d61";
		wait for Clk_period;
		Addr <=  "0001101001111";
		Trees_din <= x"00880d61";
		wait for Clk_period;
		Addr <=  "0001101010000";
		Trees_din <= x"ffd30d61";
		wait for Clk_period;
		Addr <=  "0001101010001";
		Trees_din <= x"1dffe408";
		wait for Clk_period;
		Addr <=  "0001101010010";
		Trees_din <= x"2e005404";
		wait for Clk_period;
		Addr <=  "0001101010011";
		Trees_din <= x"ff6d0d61";
		wait for Clk_period;
		Addr <=  "0001101010100";
		Trees_din <= x"fffe0d61";
		wait for Clk_period;
		Addr <=  "0001101010101";
		Trees_din <= x"2bff3204";
		wait for Clk_period;
		Addr <=  "0001101010110";
		Trees_din <= x"00520d61";
		wait for Clk_period;
		Addr <=  "0001101010111";
		Trees_din <= x"ffbd0d61";
		wait for Clk_period;
		Addr <=  "0001101011000";
		Trees_din <= x"4bff3614";
		wait for Clk_period;
		Addr <=  "0001101011001";
		Trees_din <= x"4dff5c08";
		wait for Clk_period;
		Addr <=  "0001101011010";
		Trees_din <= x"77002404";
		wait for Clk_period;
		Addr <=  "0001101011011";
		Trees_din <= x"ff6d0dd5";
		wait for Clk_period;
		Addr <=  "0001101011100";
		Trees_din <= x"00010dd5";
		wait for Clk_period;
		Addr <=  "0001101011101";
		Trees_din <= x"baffcb04";
		wait for Clk_period;
		Addr <=  "0001101011110";
		Trees_din <= x"ffb80dd5";
		wait for Clk_period;
		Addr <=  "0001101011111";
		Trees_din <= x"95ff7e04";
		wait for Clk_period;
		Addr <=  "0001101100000";
		Trees_din <= x"000b0dd5";
		wait for Clk_period;
		Addr <=  "0001101100001";
		Trees_din <= x"00570dd5";
		wait for Clk_period;
		Addr <=  "0001101100010";
		Trees_din <= x"97fec318";
		wait for Clk_period;
		Addr <=  "0001101100011";
		Trees_din <= x"1cfff210";
		wait for Clk_period;
		Addr <=  "0001101100100";
		Trees_din <= x"a3ff8e08";
		wait for Clk_period;
		Addr <=  "0001101100101";
		Trees_din <= x"35fec304";
		wait for Clk_period;
		Addr <=  "0001101100110";
		Trees_din <= x"00160dd5";
		wait for Clk_period;
		Addr <=  "0001101100111";
		Trees_din <= x"ffaf0dd5";
		wait for Clk_period;
		Addr <=  "0001101101000";
		Trees_din <= x"8cff0f04";
		wait for Clk_period;
		Addr <=  "0001101101001";
		Trees_din <= x"00590dd5";
		wait for Clk_period;
		Addr <=  "0001101101010";
		Trees_din <= x"00100dd5";
		wait for Clk_period;
		Addr <=  "0001101101011";
		Trees_din <= x"88002704";
		wait for Clk_period;
		Addr <=  "0001101101100";
		Trees_din <= x"00940dd5";
		wait for Clk_period;
		Addr <=  "0001101101101";
		Trees_din <= x"00210dd5";
		wait for Clk_period;
		Addr <=  "0001101101110";
		Trees_din <= x"48ff0e08";
		wait for Clk_period;
		Addr <=  "0001101101111";
		Trees_din <= x"11ffdb04";
		wait for Clk_period;
		Addr <=  "0001101110000";
		Trees_din <= x"00000dd5";
		wait for Clk_period;
		Addr <=  "0001101110001";
		Trees_din <= x"00590dd5";
		wait for Clk_period;
		Addr <=  "0001101110010";
		Trees_din <= x"d0ffd604";
		wait for Clk_period;
		Addr <=  "0001101110011";
		Trees_din <= x"fff50dd5";
		wait for Clk_period;
		Addr <=  "0001101110100";
		Trees_din <= x"ff870dd5";
		wait for Clk_period;
		Addr <=  "0001101110101";
		Trees_din <= x"50ff1824";
		wait for Clk_period;
		Addr <=  "0001101110110";
		Trees_din <= x"4bff5210";
		wait for Clk_period;
		Addr <=  "0001101110111";
		Trees_din <= x"a7005e08";
		wait for Clk_period;
		Addr <=  "0001101111000";
		Trees_din <= x"77ff9604";
		wait for Clk_period;
		Addr <=  "0001101111001";
		Trees_din <= x"ff8c0e39";
		wait for Clk_period;
		Addr <=  "0001101111010";
		Trees_din <= x"fff40e39";
		wait for Clk_period;
		Addr <=  "0001101111011";
		Trees_din <= x"b5feea04";
		wait for Clk_period;
		Addr <=  "0001101111100";
		Trees_din <= x"ffe10e39";
		wait for Clk_period;
		Addr <=  "0001101111101";
		Trees_din <= x"00510e39";
		wait for Clk_period;
		Addr <=  "0001101111110";
		Trees_din <= x"2effc808";
		wait for Clk_period;
		Addr <=  "0001101111111";
		Trees_din <= x"58ff3504";
		wait for Clk_period;
		Addr <=  "0001110000000";
		Trees_din <= x"ffb70e39";
		wait for Clk_period;
		Addr <=  "0001110000001";
		Trees_din <= x"00300e39";
		wait for Clk_period;
		Addr <=  "0001110000010";
		Trees_din <= x"35ff2c08";
		wait for Clk_period;
		Addr <=  "0001110000011";
		Trees_din <= x"e5fe7d04";
		wait for Clk_period;
		Addr <=  "0001110000100";
		Trees_din <= x"008b0e39";
		wait for Clk_period;
		Addr <=  "0001110000101";
		Trees_din <= x"00240e39";
		wait for Clk_period;
		Addr <=  "0001110000110";
		Trees_din <= x"00170e39";
		wait for Clk_period;
		Addr <=  "0001110000111";
		Trees_din <= x"2dffa108";
		wait for Clk_period;
		Addr <=  "0001110001000";
		Trees_din <= x"e7fee904";
		wait for Clk_period;
		Addr <=  "0001110001001";
		Trees_din <= x"ffd70e39";
		wait for Clk_period;
		Addr <=  "0001110001010";
		Trees_din <= x"ff6f0e39";
		wait for Clk_period;
		Addr <=  "0001110001011";
		Trees_din <= x"1cffde04";
		wait for Clk_period;
		Addr <=  "0001110001100";
		Trees_din <= x"ffba0e39";
		wait for Clk_period;
		Addr <=  "0001110001101";
		Trees_din <= x"00430e39";
		wait for Clk_period;
		Addr <=  "0001110001110";
		Trees_din <= x"2dff7114";
		wait for Clk_period;
		Addr <=  "0001110001111";
		Trees_din <= x"7cff070c";
		wait for Clk_period;
		Addr <=  "0001110010000";
		Trees_din <= x"2effd104";
		wait for Clk_period;
		Addr <=  "0001110010001";
		Trees_din <= x"ffaa0e95";
		wait for Clk_period;
		Addr <=  "0001110010010";
		Trees_din <= x"d6009e04";
		wait for Clk_period;
		Addr <=  "0001110010011";
		Trees_din <= x"ffed0e95";
		wait for Clk_period;
		Addr <=  "0001110010100";
		Trees_din <= x"006f0e95";
		wait for Clk_period;
		Addr <=  "0001110010101";
		Trees_din <= x"61fea404";
		wait for Clk_period;
		Addr <=  "0001110010110";
		Trees_din <= x"ffdd0e95";
		wait for Clk_period;
		Addr <=  "0001110010111";
		Trees_din <= x"ff720e95";
		wait for Clk_period;
		Addr <=  "0001110011000";
		Trees_din <= x"f4ff5f10";
		wait for Clk_period;
		Addr <=  "0001110011001";
		Trees_din <= x"1cffff08";
		wait for Clk_period;
		Addr <=  "0001110011010";
		Trees_din <= x"80fff204";
		wait for Clk_period;
		Addr <=  "0001110011011";
		Trees_din <= x"ff970e95";
		wait for Clk_period;
		Addr <=  "0001110011100";
		Trees_din <= x"00060e95";
		wait for Clk_period;
		Addr <=  "0001110011101";
		Trees_din <= x"eeff8b04";
		wait for Clk_period;
		Addr <=  "0001110011110";
		Trees_din <= x"00510e95";
		wait for Clk_period;
		Addr <=  "0001110011111";
		Trees_din <= x"00070e95";
		wait for Clk_period;
		Addr <=  "0001110100000";
		Trees_din <= x"4bfefe04";
		wait for Clk_period;
		Addr <=  "0001110100001";
		Trees_din <= x"fffb0e95";
		wait for Clk_period;
		Addr <=  "0001110100010";
		Trees_din <= x"98ff1804";
		wait for Clk_period;
		Addr <=  "0001110100011";
		Trees_din <= x"00790e95";
		wait for Clk_period;
		Addr <=  "0001110100100";
		Trees_din <= x"00110e95";
		wait for Clk_period;
		Addr <=  "0001110100101";
		Trees_din <= x"50ff181c";
		wait for Clk_period;
		Addr <=  "0001110100110";
		Trees_din <= x"54006a18";
		wait for Clk_period;
		Addr <=  "0001110100111";
		Trees_din <= x"2effb708";
		wait for Clk_period;
		Addr <=  "0001110101000";
		Trees_din <= x"f4ff4204";
		wait for Clk_period;
		Addr <=  "0001110101001";
		Trees_din <= x"ffac0ee9";
		wait for Clk_period;
		Addr <=  "0001110101010";
		Trees_din <= x"00210ee9";
		wait for Clk_period;
		Addr <=  "0001110101011";
		Trees_din <= x"daffa004";
		wait for Clk_period;
		Addr <=  "0001110101100";
		Trees_din <= x"ffe40ee9";
		wait for Clk_period;
		Addr <=  "0001110101101";
		Trees_din <= x"e5fe9408";
		wait for Clk_period;
		Addr <=  "0001110101110";
		Trees_din <= x"a0fe9904";
		wait for Clk_period;
		Addr <=  "0001110101111";
		Trees_din <= x"00180ee9";
		wait for Clk_period;
		Addr <=  "0001110110000";
		Trees_din <= x"00810ee9";
		wait for Clk_period;
		Addr <=  "0001110110001";
		Trees_din <= x"000a0ee9";
		wait for Clk_period;
		Addr <=  "0001110110010";
		Trees_din <= x"ffa40ee9";
		wait for Clk_period;
		Addr <=  "0001110110011";
		Trees_din <= x"17ff4e08";
		wait for Clk_period;
		Addr <=  "0001110110100";
		Trees_din <= x"97febd04";
		wait for Clk_period;
		Addr <=  "0001110110101";
		Trees_din <= x"004c0ee9";
		wait for Clk_period;
		Addr <=  "0001110110110";
		Trees_din <= x"ffd20ee9";
		wait for Clk_period;
		Addr <=  "0001110110111";
		Trees_din <= x"2dffdd04";
		wait for Clk_period;
		Addr <=  "0001110111000";
		Trees_din <= x"ff730ee9";
		wait for Clk_period;
		Addr <=  "0001110111001";
		Trees_din <= x"fff90ee9";
		wait for Clk_period;
		Addr <=  "0001110111010";
		Trees_din <= x"1cffd914";
		wait for Clk_period;
		Addr <=  "0001110111011";
		Trees_din <= x"48fea308";
		wait for Clk_period;
		Addr <=  "0001110111100";
		Trees_din <= x"2affc504";
		wait for Clk_period;
		Addr <=  "0001110111101";
		Trees_din <= x"00500f35";
		wait for Clk_period;
		Addr <=  "0001110111110";
		Trees_din <= x"fff30f35";
		wait for Clk_period;
		Addr <=  "0001110111111";
		Trees_din <= x"2dff9e04";
		wait for Clk_period;
		Addr <=  "0001111000000";
		Trees_din <= x"ff750f35";
		wait for Clk_period;
		Addr <=  "0001111000001";
		Trees_din <= x"bafffd04";
		wait for Clk_period;
		Addr <=  "0001111000010";
		Trees_din <= x"ffbf0f35";
		wait for Clk_period;
		Addr <=  "0001111000011";
		Trees_din <= x"001d0f35";
		wait for Clk_period;
		Addr <=  "0001111000100";
		Trees_din <= x"17ffcc10";
		wait for Clk_period;
		Addr <=  "0001111000101";
		Trees_din <= x"02fee504";
		wait for Clk_period;
		Addr <=  "0001111000110";
		Trees_din <= x"ffe90f35";
		wait for Clk_period;
		Addr <=  "0001111000111";
		Trees_din <= x"e3febf08";
		wait for Clk_period;
		Addr <=  "0001111001000";
		Trees_din <= x"1f002904";
		wait for Clk_period;
		Addr <=  "0001111001001";
		Trees_din <= x"007b0f35";
		wait for Clk_period;
		Addr <=  "0001111001010";
		Trees_din <= x"00210f35";
		wait for Clk_period;
		Addr <=  "0001111001011";
		Trees_din <= x"00100f35";
		wait for Clk_period;
		Addr <=  "0001111001100";
		Trees_din <= x"ffbb0f35";
		wait for Clk_period;
		Addr <=  "0001111001101";
		Trees_din <= x"a700080c";
		wait for Clk_period;
		Addr <=  "0001111001110";
		Trees_din <= x"02ffd908";
		wait for Clk_period;
		Addr <=  "0001111001111";
		Trees_din <= x"17ff3b04";
		wait for Clk_period;
		Addr <=  "0001111010000";
		Trees_din <= x"00010f81";
		wait for Clk_period;
		Addr <=  "0001111010001";
		Trees_din <= x"ff750f81";
		wait for Clk_period;
		Addr <=  "0001111010010";
		Trees_din <= x"00370f81";
		wait for Clk_period;
		Addr <=  "0001111010011";
		Trees_din <= x"4bff0508";
		wait for Clk_period;
		Addr <=  "0001111010100";
		Trees_din <= x"d4ffa804";
		wait for Clk_period;
		Addr <=  "0001111010101";
		Trees_din <= x"ff9e0f81";
		wait for Clk_period;
		Addr <=  "0001111010110";
		Trees_din <= x"00240f81";
		wait for Clk_period;
		Addr <=  "0001111010111";
		Trees_din <= x"f4fef204";
		wait for Clk_period;
		Addr <=  "0001111011000";
		Trees_din <= x"ffeb0f81";
		wait for Clk_period;
		Addr <=  "0001111011001";
		Trees_din <= x"01fde804";
		wait for Clk_period;
		Addr <=  "0001111011010";
		Trees_din <= x"fffc0f81";
		wait for Clk_period;
		Addr <=  "0001111011011";
		Trees_din <= x"1dff6f04";
		wait for Clk_period;
		Addr <=  "0001111011100";
		Trees_din <= x"00080f81";
		wait for Clk_period;
		Addr <=  "0001111011101";
		Trees_din <= x"35ff1404";
		wait for Clk_period;
		Addr <=  "0001111011110";
		Trees_din <= x"00770f81";
		wait for Clk_period;
		Addr <=  "0001111011111";
		Trees_din <= x"00200f81";
		wait for Clk_period;
		Addr <=  "0001111100000";
		Trees_din <= x"4bff350c";
		wait for Clk_period;
		Addr <=  "0001111100001";
		Trees_din <= x"4dff5c08";
		wait for Clk_period;
		Addr <=  "0001111100010";
		Trees_din <= x"1dffa404";
		wait for Clk_period;
		Addr <=  "0001111100011";
		Trees_din <= x"ff770fbd";
		wait for Clk_period;
		Addr <=  "0001111100100";
		Trees_din <= x"ffdc0fbd";
		wait for Clk_period;
		Addr <=  "0001111100101";
		Trees_din <= x"00150fbd";
		wait for Clk_period;
		Addr <=  "0001111100110";
		Trees_din <= x"97fecc0c";
		wait for Clk_period;
		Addr <=  "0001111100111";
		Trees_din <= x"84001008";
		wait for Clk_period;
		Addr <=  "0001111101000";
		Trees_din <= x"2a002304";
		wait for Clk_period;
		Addr <=  "0001111101001";
		Trees_din <= x"00740fbd";
		wait for Clk_period;
		Addr <=  "0001111101010";
		Trees_din <= x"00120fbd";
		wait for Clk_period;
		Addr <=  "0001111101011";
		Trees_din <= x"fff90fbd";
		wait for Clk_period;
		Addr <=  "0001111101100";
		Trees_din <= x"7cff0204";
		wait for Clk_period;
		Addr <=  "0001111101101";
		Trees_din <= x"00310fbd";
		wait for Clk_period;
		Addr <=  "0001111101110";
		Trees_din <= x"ff9e0fbd";
		wait for Clk_period;
		Addr <=  "0001111101111";
		Trees_din <= x"50ff1818";
		wait for Clk_period;
		Addr <=  "0001111110000";
		Trees_din <= x"54006a14";
		wait for Clk_period;
		Addr <=  "0001111110001";
		Trees_din <= x"2effb708";
		wait for Clk_period;
		Addr <=  "0001111110010";
		Trees_din <= x"acffe304";
		wait for Clk_period;
		Addr <=  "0001111110011";
		Trees_din <= x"00261001";
		wait for Clk_period;
		Addr <=  "0001111110100";
		Trees_din <= x"ffc11001";
		wait for Clk_period;
		Addr <=  "0001111110101";
		Trees_din <= x"eaff4604";
		wait for Clk_period;
		Addr <=  "0001111110110";
		Trees_din <= x"fff61001";
		wait for Clk_period;
		Addr <=  "0001111110111";
		Trees_din <= x"e5fe9104";
		wait for Clk_period;
		Addr <=  "0001111111000";
		Trees_din <= x"006a1001";
		wait for Clk_period;
		Addr <=  "0001111111001";
		Trees_din <= x"000c1001";
		wait for Clk_period;
		Addr <=  "0001111111010";
		Trees_din <= x"ffb71001";
		wait for Clk_period;
		Addr <=  "0001111111011";
		Trees_din <= x"1dffe408";
		wait for Clk_period;
		Addr <=  "0001111111100";
		Trees_din <= x"fcffa204";
		wait for Clk_period;
		Addr <=  "0001111111101";
		Trees_din <= x"ff791001";
		wait for Clk_period;
		Addr <=  "0001111111110";
		Trees_din <= x"fff01001";
		wait for Clk_period;
		Addr <=  "0001111111111";
		Trees_din <= x"001b1001";
		wait for Clk_period;
		Addr <=  "0010000000000";
		Trees_din <= x"78ffe710";
		wait for Clk_period;
		Addr <=  "0010000000001";
		Trees_din <= x"1c002d0c";
		wait for Clk_period;
		Addr <=  "0010000000010";
		Trees_din <= x"06fe9904";
		wait for Clk_period;
		Addr <=  "0010000000011";
		Trees_din <= x"0001103d";
		wait for Clk_period;
		Addr <=  "0010000000100";
		Trees_din <= x"e7ff0d04";
		wait for Clk_period;
		Addr <=  "0010000000101";
		Trees_din <= x"ffd5103d";
		wait for Clk_period;
		Addr <=  "0010000000110";
		Trees_din <= x"ff7b103d";
		wait for Clk_period;
		Addr <=  "0010000000111";
		Trees_din <= x"0030103d";
		wait for Clk_period;
		Addr <=  "0010000001000";
		Trees_din <= x"d0001308";
		wait for Clk_period;
		Addr <=  "0010000001001";
		Trees_din <= x"e1ffa504";
		wait for Clk_period;
		Addr <=  "0010000001010";
		Trees_din <= x"000e103d";
		wait for Clk_period;
		Addr <=  "0010000001011";
		Trees_din <= x"0064103d";
		wait for Clk_period;
		Addr <=  "0010000001100";
		Trees_din <= x"2bfe5a04";
		wait for Clk_period;
		Addr <=  "0010000001101";
		Trees_din <= x"0032103d";
		wait for Clk_period;
		Addr <=  "0010000001110";
		Trees_din <= x"ffbb103d";
		wait for Clk_period;
		Addr <=  "0010000001111";
		Trees_din <= x"a700080c";
		wait for Clk_period;
		Addr <=  "0010000010000";
		Trees_din <= x"4bff5504";
		wait for Clk_period;
		Addr <=  "0010000010001";
		Trees_din <= x"ff831081";
		wait for Clk_period;
		Addr <=  "0010000010010";
		Trees_din <= x"bffefe04";
		wait for Clk_period;
		Addr <=  "0010000010011";
		Trees_din <= x"003c1081";
		wait for Clk_period;
		Addr <=  "0010000010100";
		Trees_din <= x"ffbf1081";
		wait for Clk_period;
		Addr <=  "0010000010101";
		Trees_din <= x"1cffff10";
		wait for Clk_period;
		Addr <=  "0010000010110";
		Trees_din <= x"80ffde08";
		wait for Clk_period;
		Addr <=  "0010000010111";
		Trees_din <= x"e7feff04";
		wait for Clk_period;
		Addr <=  "0010000011000";
		Trees_din <= x"000c1081";
		wait for Clk_period;
		Addr <=  "0010000011001";
		Trees_din <= x"ffac1081";
		wait for Clk_period;
		Addr <=  "0010000011010";
		Trees_din <= x"22ff1404";
		wait for Clk_period;
		Addr <=  "0010000011011";
		Trees_din <= x"004e1081";
		wait for Clk_period;
		Addr <=  "0010000011100";
		Trees_din <= x"fff51081";
		wait for Clk_period;
		Addr <=  "0010000011101";
		Trees_din <= x"1dffce04";
		wait for Clk_period;
		Addr <=  "0010000011110";
		Trees_din <= x"00151081";
		wait for Clk_period;
		Addr <=  "0010000011111";
		Trees_din <= x"00641081";
		wait for Clk_period;
		Addr <=  "0010000100000";
		Trees_din <= x"e7ff1a0c";
		wait for Clk_period;
		Addr <=  "0010000100001";
		Trees_din <= x"17ffd908";
		wait for Clk_period;
		Addr <=  "0010000100010";
		Trees_din <= x"8cff7304";
		wait for Clk_period;
		Addr <=  "0010000100011";
		Trees_din <= x"006510ad";
		wait for Clk_period;
		Addr <=  "0010000100100";
		Trees_din <= x"000e10ad";
		wait for Clk_period;
		Addr <=  "0010000100101";
		Trees_din <= x"ffd810ad";
		wait for Clk_period;
		Addr <=  "0010000100110";
		Trees_din <= x"94009c08";
		wait for Clk_period;
		Addr <=  "0010000100111";
		Trees_din <= x"4bffac04";
		wait for Clk_period;
		Addr <=  "0010000101000";
		Trees_din <= x"ff8410ad";
		wait for Clk_period;
		Addr <=  "0010000101001";
		Trees_din <= x"000a10ad";
		wait for Clk_period;
		Addr <=  "0010000101010";
		Trees_din <= x"002010ad";
		wait for Clk_period;
		Addr <=  "0010000101011";
		Trees_din <= x"a700080c";
		wait for Clk_period;
		Addr <=  "0010000101100";
		Trees_din <= x"1cffd904";
		wait for Clk_period;
		Addr <=  "0010000101101";
		Trees_din <= x"ff8a10e1";
		wait for Clk_period;
		Addr <=  "0010000101110";
		Trees_din <= x"bffefe04";
		wait for Clk_period;
		Addr <=  "0010000101111";
		Trees_din <= x"003110e1";
		wait for Clk_period;
		Addr <=  "0010000110000";
		Trees_din <= x"ffc710e1";
		wait for Clk_period;
		Addr <=  "0010000110001";
		Trees_din <= x"d0006c0c";
		wait for Clk_period;
		Addr <=  "0010000110010";
		Trees_din <= x"4dfeab04";
		wait for Clk_period;
		Addr <=  "0010000110011";
		Trees_din <= x"fff010e1";
		wait for Clk_period;
		Addr <=  "0010000110100";
		Trees_din <= x"b8ff4c04";
		wait for Clk_period;
		Addr <=  "0010000110101";
		Trees_din <= x"005b10e1";
		wait for Clk_period;
		Addr <=  "0010000110110";
		Trees_din <= x"000810e1";
		wait for Clk_period;
		Addr <=  "0010000110111";
		Trees_din <= x"ffd910e1";
		wait for Clk_period;
		Addr <=  "0010000111000";
		Trees_din <= x"50ff1814";
		wait for Clk_period;
		Addr <=  "0010000111001";
		Trees_din <= x"80ff8a04";
		wait for Clk_period;
		Addr <=  "0010000111010";
		Trees_din <= x"ffd6111d";
		wait for Clk_period;
		Addr <=  "0010000111011";
		Trees_din <= x"cafe3404";
		wait for Clk_period;
		Addr <=  "0010000111100";
		Trees_din <= x"ffe9111d";
		wait for Clk_period;
		Addr <=  "0010000111101";
		Trees_din <= x"88001e08";
		wait for Clk_period;
		Addr <=  "0010000111110";
		Trees_din <= x"1cffab04";
		wait for Clk_period;
		Addr <=  "0010000111111";
		Trees_din <= x"001f111d";
		wait for Clk_period;
		Addr <=  "0010001000000";
		Trees_din <= x"006a111d";
		wait for Clk_period;
		Addr <=  "0010001000001";
		Trees_din <= x"0005111d";
		wait for Clk_period;
		Addr <=  "0010001000010";
		Trees_din <= x"1dffe408";
		wait for Clk_period;
		Addr <=  "0010001000011";
		Trees_din <= x"e4fe1904";
		wait for Clk_period;
		Addr <=  "0010001000100";
		Trees_din <= x"ffe8111d";
		wait for Clk_period;
		Addr <=  "0010001000101";
		Trees_din <= x"ff86111d";
		wait for Clk_period;
		Addr <=  "0010001000110";
		Trees_din <= x"0018111d";
		wait for Clk_period;
		Addr <=  "0010001000111";
		Trees_din <= x"48ff1208";
		wait for Clk_period;
		Addr <=  "0010001001000";
		Trees_din <= x"2a000f04";
		wait for Clk_period;
		Addr <=  "0010001001001";
		Trees_din <= x"00561149";
		wait for Clk_period;
		Addr <=  "0010001001010";
		Trees_din <= x"ffee1149";
		wait for Clk_period;
		Addr <=  "0010001001011";
		Trees_din <= x"2dff9008";
		wait for Clk_period;
		Addr <=  "0010001001100";
		Trees_din <= x"e7ff1504";
		wait for Clk_period;
		Addr <=  "0010001001101";
		Trees_din <= x"fff31149";
		wait for Clk_period;
		Addr <=  "0010001001110";
		Trees_din <= x"ff861149";
		wait for Clk_period;
		Addr <=  "0010001001111";
		Trees_din <= x"9bff5804";
		wait for Clk_period;
		Addr <=  "0010001010000";
		Trees_din <= x"ffd91149";
		wait for Clk_period;
		Addr <=  "0010001010001";
		Trees_din <= x"00381149";
		wait for Clk_period;
		Addr <=  "0010001010010";
		Trees_din <= x"4bff3508";
		wait for Clk_period;
		Addr <=  "0010001010011";
		Trees_din <= x"4dff5c04";
		wait for Clk_period;
		Addr <=  "0010001010100";
		Trees_din <= x"ff96117d";
		wait for Clk_period;
		Addr <=  "0010001010101";
		Trees_din <= x"0011117d";
		wait for Clk_period;
		Addr <=  "0010001010110";
		Trees_din <= x"f4fef104";
		wait for Clk_period;
		Addr <=  "0010001010111";
		Trees_din <= x"ffd1117d";
		wait for Clk_period;
		Addr <=  "0010001011000";
		Trees_din <= x"bfff2208";
		wait for Clk_period;
		Addr <=  "0010001011001";
		Trees_din <= x"1cffe204";
		wait for Clk_period;
		Addr <=  "0010001011010";
		Trees_din <= x"0016117d";
		wait for Clk_period;
		Addr <=  "0010001011011";
		Trees_din <= x"0062117d";
		wait for Clk_period;
		Addr <=  "0010001011100";
		Trees_din <= x"1dffc104";
		wait for Clk_period;
		Addr <=  "0010001011101";
		Trees_din <= x"ffe2117d";
		wait for Clk_period;
		Addr <=  "0010001011110";
		Trees_din <= x"0020117d";
		wait for Clk_period;
		Addr <=  "0010001011111";
		Trees_din <= x"d000230c";
		wait for Clk_period;
		Addr <=  "0010001100000";
		Trees_din <= x"71ff0908";
		wait for Clk_period;
		Addr <=  "0010001100001";
		Trees_din <= x"2a000f04";
		wait for Clk_period;
		Addr <=  "0010001100010";
		Trees_din <= x"005411a9";
		wait for Clk_period;
		Addr <=  "0010001100011";
		Trees_din <= x"000411a9";
		wait for Clk_period;
		Addr <=  "0010001100100";
		Trees_din <= x"ffe011a9";
		wait for Clk_period;
		Addr <=  "0010001100101";
		Trees_din <= x"4c002308";
		wait for Clk_period;
		Addr <=  "0010001100110";
		Trees_din <= x"4dff0b04";
		wait for Clk_period;
		Addr <=  "0010001100111";
		Trees_din <= x"ff9111a9";
		wait for Clk_period;
		Addr <=  "0010001101000";
		Trees_din <= x"fff211a9";
		wait for Clk_period;
		Addr <=  "0010001101001";
		Trees_din <= x"001a11a9";
		wait for Clk_period;
		Addr <=  "0010001101010";
		Trees_din <= x"48ff120c";
		wait for Clk_period;
		Addr <=  "0010001101011";
		Trees_din <= x"47000508";
		wait for Clk_period;
		Addr <=  "0010001101100";
		Trees_din <= x"83fef904";
		wait for Clk_period;
		Addr <=  "0010001101101";
		Trees_din <= x"005811d5";
		wait for Clk_period;
		Addr <=  "0010001101110";
		Trees_din <= x"001511d5";
		wait for Clk_period;
		Addr <=  "0010001101111";
		Trees_din <= x"ffe611d5";
		wait for Clk_period;
		Addr <=  "0010001110000";
		Trees_din <= x"97fec908";
		wait for Clk_period;
		Addr <=  "0010001110001";
		Trees_din <= x"1cfff204";
		wait for Clk_period;
		Addr <=  "0010001110010";
		Trees_din <= x"ffdb11d5";
		wait for Clk_period;
		Addr <=  "0010001110011";
		Trees_din <= x"003a11d5";
		wait for Clk_period;
		Addr <=  "0010001110100";
		Trees_din <= x"ff9c11d5";
		wait for Clk_period;
		Addr <=  "0010001110101";
		Trees_din <= x"78ffe70c";
		wait for Clk_period;
		Addr <=  "0010001110110";
		Trees_din <= x"06fea204";
		wait for Clk_period;
		Addr <=  "0010001110111";
		Trees_din <= x"00201201";
		wait for Clk_period;
		Addr <=  "0010001111000";
		Trees_din <= x"2dff7604";
		wait for Clk_period;
		Addr <=  "0010001111001";
		Trees_din <= x"ff931201";
		wait for Clk_period;
		Addr <=  "0010001111010";
		Trees_din <= x"ffef1201";
		wait for Clk_period;
		Addr <=  "0010001111011";
		Trees_din <= x"6bff0d08";
		wait for Clk_period;
		Addr <=  "0010001111100";
		Trees_din <= x"d0004104";
		wait for Clk_period;
		Addr <=  "0010001111101";
		Trees_din <= x"00531201";
		wait for Clk_period;
		Addr <=  "0010001111110";
		Trees_din <= x"fff61201";
		wait for Clk_period;
		Addr <=  "0010001111111";
		Trees_din <= x"ffe81201";
		wait for Clk_period;
		Addr <=  "0010010000000";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  7
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"1f011f80";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"ab008e40";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"20004020";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"8c00b010";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"75004808";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"f0fffe04";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"ff82014d";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"000a014d";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"d0014f04";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"ffbe014d";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"0117014d";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"31ffda08";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"83ff2e04";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"000f014d";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"030a014d";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"7cff2204";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"0114014d";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"ff79014d";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"01feaa10";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"c9ffe408";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"3d005d04";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"ffe1014d";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"01b7014d";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"66ffb104";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"fff8014d";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"0215014d";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"2b003008";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"ba003004";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"ff81014d";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"00cd014d";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"21000904";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"022f014d";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"ff96014d";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"31000420";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"2fffe610";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"5a004308";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"af002104";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"0007014d";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"015e014d";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"11ffd504";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"ff9d014d";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"00cc014d";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"aefee008";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"21001904";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"ff93014d";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"00ed014d";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"65fe7d04";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"ff66014d";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"014d014d";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"4bfee310";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"2fffa108";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"6aff2704";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"01f5014d";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"ffaa014d";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"b9fee204";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"ffea014d";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"0206014d";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"eeffab08";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"c2ff8704";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"ffc1014d";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"0192014d";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"4effbd04";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"012c014d";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"031d014d";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"01fe8014";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"bdffca0c";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"d8009c08";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"80fef804";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"00ca014d";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"041b014d";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"0021014d";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"c2ffa704";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"ff81014d";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"01f5014d";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"faff8408";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"faff0504";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"015c014d";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"ff65014d";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"c5ff3504";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"030a014d";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"75005504";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"ff73014d";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"01f5014d";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"1f00e77c";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"ab00ef40";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"1fffcd20";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"73ffea10";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"99006708";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"07013e04";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"ff8f0299";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"00d80299";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"1dff9904";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"ff850299";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"01fd0299";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"b1ff0808";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"c7ff6104";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"ffdf0299";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"00ee0299";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"75006604";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"ff820299";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"001a0299";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"00ff6e10";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"a4ff1408";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"6e006204";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"01610299";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"ff990299";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"1afe9204";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"00200299";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"ff9d0299";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"84ff8a08";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"1b007d04";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"ffcb0299";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"00f70299";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"59ff7a04";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"00e40299";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"000e0299";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"feff8a1c";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"a1fec410";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"89ffdc08";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"b7fff504";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"ff660299";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"00ed0299";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"62ff3a04";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"002d0299";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"02610299";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"adfefc04";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"015d0299";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"5affaf04";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"00d70299";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"ff6a0299";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"aefedf10";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"54001808";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"00ff5b04";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"ff840299";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"01b70299";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"d2fe4704";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"00ac0299";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"ff5c0299";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"03ff7b08";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"3d000304";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"ffa20299";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"01610299";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"43ffab04";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"01ca0299";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"fff70299";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"66ff770c";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"1dfea308";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"c9ffb804";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"00d70299";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"00390299";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"ff630299";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"00ff2208";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"2efff104";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"ff6a0299";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"00f90299";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"91fff910";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"f8ffe108";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"12ff9b04";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"003b0299";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"ff870299";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"e7ffd604";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"01b40299";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"fff40299";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"b2ff5b04";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"00380299";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"ff800299";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"01fe7b7c";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"20fff740";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"ab00ac20";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"8dff1510";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"5400a108";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"8c004504";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"ff8a0485";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"003e0485";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"14feef04";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"ffb00485";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"01170485";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"b3ff1008";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"ddff8504";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"ff760485";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"003b0485";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"4aff8004";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"020b0485";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"ff990485";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"30ffff10";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"11ffb308";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"7aff1f04";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"00e40485";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"ff990485";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"0a007804";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"017e0485";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"ffc70485";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"8cff4208";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"dc008f04";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"ff670485";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"00b70485";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"c7fe9004";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"004d0485";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"01b00485";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"4dfef820";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"d8002810";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"e6ffa308";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"62ff6304";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"01590485";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"ffb30485";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"0800aa04";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"ff620485";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"005f0485";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"4efe5008";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"e1005a04";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"ff700485";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"00a40485";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"64ff6004";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"018a0485";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"00880485";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"3eff460c";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"71ff6808";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"9fffa804";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"ff800485";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"00c10485";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"01ef0485";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"90ff0408";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"8dfdf804";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"01500485";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"ff9c0485";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"3bfe0c04";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"00290485";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"ff5c0485";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"10ffe83c";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"b6ff721c";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"26010910";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"d2ff7508";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"c3ff1c04";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"00430485";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"ff810485";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"47fff604";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"ff940485";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"01500485";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"73000204";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"01e30485";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"66001b04";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"ff9a0485";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"00340485";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"b3ff7110";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"9cffd108";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"00ff9d04";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"ff7b0485";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"00020485";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"53ff2a04";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"01420485";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"ffdb0485";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"29ff7b08";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"13004004";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"00f00485";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"ff780485";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"deffd304";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"02100485";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"00650485";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"69fed820";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"1effb710";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"2dfeb108";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"5bff7a04";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"00410485";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"021f0485";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"c2ffd204";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"ff830485";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"009b0485";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"60ff5a08";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"bcfef004";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"01250485";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"ff700485";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"b5fef204";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"021d0485";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"00310485";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"a9fede10";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"3eff9708";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"3f004c04";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"ff880485";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"014b0485";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"11ff6704";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"02ad0485";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"00370485";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"ab00b308";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"2e004204";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"ffa30485";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"00900485";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"5cff7804";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"01470485";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"00080485";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"01fe7b70";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"1f002438";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"28ff3920";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"1300ec10";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"8cff7908";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"5ffee204";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"00330641";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"ff740641";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"4effd104";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"00020641";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"00ee0641";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"6c004e08";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"87ffee04";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"ff6d0641";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"009a0641";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"b6ff6204";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"01670641";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"ffa20641";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"d8001b0c";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"2dfde804";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"00c60641";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"40ff9104";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"009f0641";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"ff5e0641";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"58ff6e08";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"49ffa304";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"01430641";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"00600641";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"ff6d0641";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"83ff3720";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"3bff1a10";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"7efe6c08";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"1dffa104";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"018d0641";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"ff9e0641";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"a6ff4304";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"00e60641";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"ff6a0641";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"34004408";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"e3fedc04";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"ff8c0641";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"00890641";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"83ff0a04";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"013b0641";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"ff920641";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"6a000210";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"56ff7e08";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"39006c04";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"01150641";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"ff8b0641";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"04009c04";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"ffa30641";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"01400641";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"84002204";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"ff680641";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"00d10641";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"0b005b40";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"75005420";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"89009e10";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"2f000208";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"27ff0404";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"00390641";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"ffa00641";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"c0ff5104";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"00ee0641";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"ffc00641";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"66ffe108";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"35fec604";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"ff800641";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"011d0641";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"82ffca04";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"ff660641";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"00b90641";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"b6ffbe10";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"55001e08";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"ea001504";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"ff8e0641";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"00a80641";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"79ff6104";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"005f0641";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"ffa90641";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"ecffe708";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"dc006f04";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"ff6d0641";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"00a00641";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"b2ff9104";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"ff840641";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"018a0641";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"ab00731c";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"a4ff510c";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"f0ff2e04";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"ff710641";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"10004604";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"00190641";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"01c60641";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"94ff5308";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"0a002004";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"01d30641";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"ff930641";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"98ffab04";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"ff710641";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"009a0641";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"31ff5704";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"ff700641";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"cb002d08";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"84ff6004";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"ff8e0641";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"017f0641";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"12ffab04";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"00fb0641";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"ff830641";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"01fe7e64";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"20fff740";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"11ff7420";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"a0ff6810";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"1afe9608";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"c3ffd104";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"00a707fd";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"ff9107fd";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"43fea304";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"006d07fd";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"ff8d07fd";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"1300a308";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"07008604";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"ff7907fd";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"003407fd";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"ab004d04";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"000507fd";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"01a807fd";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"45fe7910";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"15ff3108";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"effeed04";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"01aa07fd";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"ffe007fd";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"d000e904";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"ff6b07fd";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"004607fd";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"ebff1208";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"f8002104";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"ff9e07fd";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"009807fd";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"9a001704";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"015307fd";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"ff8207fd";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"6a001e20";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"44ff9310";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"20005e08";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"e2fe4604";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"003207fd";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"ff5d07fd";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"36ff2004";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"ff9a07fd";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"00c107fd";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"b5ff0b08";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"64ff5a04";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"00a007fd";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"ffdd07fd";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"78ffcd04";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"015c07fd";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"003207fd";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"ff6f07fd";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"10ffe83c";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"a8ff2b1c";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"1afeea0c";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"20ff3c04";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"ff6b07fd";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"77feb904";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"ffa007fd";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"00a607fd";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"b8001708";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"8800ba04";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"ff7f07fd";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"009a07fd";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"e3fe6e04";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"020c07fd";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"ff8e07fd";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"66004d10";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"c0fff608";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"2ffff104";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"ff8c07fd";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"001707fd";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"5dff4a04";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"01d007fd";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"ffd807fd";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"13008808";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"9afffc04";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"01a007fd";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"ff8c07fd";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"58fe6b04";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"00b407fd";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"ff6507fd";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"6bfe9b20";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"64fec710";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"a1feb108";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"9eff7f04";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"01ee07fd";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"002707fd";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"73000f04";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"ff6c07fd";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"008107fd";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"d1feff08";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"45ff0c04";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"011e07fd";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"ff8807fd";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"cf00dc04";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"ff7f07fd";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"009607fd";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"69ff0d10";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"e9ff4508";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"66ff7704";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"ffc207fd";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"00f807fd";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"28fea904";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"00d007fd";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"ff6c07fd";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"d4fef508";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"83ff9304";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"016207fd";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"ff8607fd";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"d9ffe604";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"ffc807fd";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"006307fd";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"8cffe07c";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"c2ffc240";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"ab00cd20";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"20003210";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"b5005308";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"24008b04";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"ffa609c9";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"007e09c9";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"0dff3e04";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"ffa209c9";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"01e709c9";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"7aff9b08";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"7aff5c04";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"ffc509c9";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"012009c9";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"11ffd304";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"ff7709c9";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"00c409c9";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"f7ff2110";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"1bffc808";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"00ffc904";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"ff9b09c9";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"010709c9";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"3fffe404";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"ff7909c9";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"010509c9";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"19feee08";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"f6fe9904";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"01c809c9";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"ffdb09c9";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"c8006f04";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"ff7209c9";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"006209c9";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"3ffffe20";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"20fff210";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"a5feab08";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"f4fef404";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"ff8209c9";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"00f609c9";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"7200af04";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"ff6a09c9";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"009d09c9";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"5fff4308";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"8dfdf904";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"00b909c9";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"ff7809c9";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"10ff2e04";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"001709c9";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"018f09c9";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"61ff7a10";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"92ff7f08";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"02fe6104";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"00da09c9";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"ffd209c9";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"12ff9e04";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"01d009c9";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"001409c9";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"e4ff3108";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"1aff2004";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"014e09c9";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"ffbb09c9";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"ff7809c9";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"6fff4130";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"4dfe5210";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"9dff3804";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"ff7b09c9";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"19ffad08";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"0cfe5904";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"003a09c9";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"013109c9";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"ff8909c9";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"5cffce10";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"f9ff2608";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"ddff5d04";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"ffaf09c9";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"00d609c9";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"66ff6204";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"ff9d09c9";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"017a09c9";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"5100b608";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"8c003504";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"ff8809c9";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"002509c9";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"a8ff9a04";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"010309c9";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"ff8409c9";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"90ff541c";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"01fde80c";
		wait for Clk_period;
		Addr <=  "0001001010111";
		Trees_din <= x"87ff2604";
		wait for Clk_period;
		Addr <=  "0001001011000";
		Trees_din <= x"ff8d09c9";
		wait for Clk_period;
		Addr <=  "0001001011001";
		Trees_din <= x"49ffec04";
		wait for Clk_period;
		Addr <=  "0001001011010";
		Trees_din <= x"006009c9";
		wait for Clk_period;
		Addr <=  "0001001011011";
		Trees_din <= x"016a09c9";
		wait for Clk_period;
		Addr <=  "0001001011100";
		Trees_din <= x"72ffc508";
		wait for Clk_period;
		Addr <=  "0001001011101";
		Trees_din <= x"b4ff2404";
		wait for Clk_period;
		Addr <=  "0001001011110";
		Trees_din <= x"00ad09c9";
		wait for Clk_period;
		Addr <=  "0001001011111";
		Trees_din <= x"ffb109c9";
		wait for Clk_period;
		Addr <=  "0001001100000";
		Trees_din <= x"9bff2104";
		wait for Clk_period;
		Addr <=  "0001001100001";
		Trees_din <= x"fff209c9";
		wait for Clk_period;
		Addr <=  "0001001100010";
		Trees_din <= x"ff7e09c9";
		wait for Clk_period;
		Addr <=  "0001001100011";
		Trees_din <= x"b0ffb710";
		wait for Clk_period;
		Addr <=  "0001001100100";
		Trees_din <= x"f0004608";
		wait for Clk_period;
		Addr <=  "0001001100101";
		Trees_din <= x"b4ff0804";
		wait for Clk_period;
		Addr <=  "0001001100110";
		Trees_din <= x"003809c9";
		wait for Clk_period;
		Addr <=  "0001001100111";
		Trees_din <= x"ffb409c9";
		wait for Clk_period;
		Addr <=  "0001001101000";
		Trees_din <= x"90fff204";
		wait for Clk_period;
		Addr <=  "0001001101001";
		Trees_din <= x"01bf09c9";
		wait for Clk_period;
		Addr <=  "0001001101010";
		Trees_din <= x"000209c9";
		wait for Clk_period;
		Addr <=  "0001001101011";
		Trees_din <= x"ab005208";
		wait for Clk_period;
		Addr <=  "0001001101100";
		Trees_din <= x"db009b04";
		wait for Clk_period;
		Addr <=  "0001001101101";
		Trees_din <= x"ffa009c9";
		wait for Clk_period;
		Addr <=  "0001001101110";
		Trees_din <= x"00d409c9";
		wait for Clk_period;
		Addr <=  "0001001101111";
		Trees_din <= x"eaff7304";
		wait for Clk_period;
		Addr <=  "0001001110000";
		Trees_din <= x"000f09c9";
		wait for Clk_period;
		Addr <=  "0001001110001";
		Trees_din <= x"013d09c9";
		wait for Clk_period;
		Addr <=  "0001001110010";
		Trees_din <= x"89008a74";
		wait for Clk_period;
		Addr <=  "0001001110011";
		Trees_din <= x"ab008e34";
		wait for Clk_period;
		Addr <=  "0001001110100";
		Trees_din <= x"f0004620";
		wait for Clk_period;
		Addr <=  "0001001110101";
		Trees_din <= x"09ffdb10";
		wait for Clk_period;
		Addr <=  "0001001110110";
		Trees_din <= x"d5001508";
		wait for Clk_period;
		Addr <=  "0001001110111";
		Trees_din <= x"2700b204";
		wait for Clk_period;
		Addr <=  "0001001111000";
		Trees_din <= x"ff8f0b65";
		wait for Clk_period;
		Addr <=  "0001001111001";
		Trees_din <= x"007a0b65";
		wait for Clk_period;
		Addr <=  "0001001111010";
		Trees_din <= x"f8005d04";
		wait for Clk_period;
		Addr <=  "0001001111011";
		Trees_din <= x"ffb90b65";
		wait for Clk_period;
		Addr <=  "0001001111100";
		Trees_din <= x"00560b65";
		wait for Clk_period;
		Addr <=  "0001001111101";
		Trees_din <= x"30ff6b08";
		wait for Clk_period;
		Addr <=  "0001001111110";
		Trees_din <= x"25009304";
		wait for Clk_period;
		Addr <=  "0001001111111";
		Trees_din <= x"ff620b65";
		wait for Clk_period;
		Addr <=  "0001010000000";
		Trees_din <= x"00440b65";
		wait for Clk_period;
		Addr <=  "0001010000001";
		Trees_din <= x"a1fefc04";
		wait for Clk_period;
		Addr <=  "0001010000010";
		Trees_din <= x"ffc70b65";
		wait for Clk_period;
		Addr <=  "0001010000011";
		Trees_din <= x"004e0b65";
		wait for Clk_period;
		Addr <=  "0001010000100";
		Trees_din <= x"bcff8510";
		wait for Clk_period;
		Addr <=  "0001010000101";
		Trees_din <= x"6fffa608";
		wait for Clk_period;
		Addr <=  "0001010000110";
		Trees_din <= x"4cff2804";
		wait for Clk_period;
		Addr <=  "0001010000111";
		Trees_din <= x"00d30b65";
		wait for Clk_period;
		Addr <=  "0001010001000";
		Trees_din <= x"ff8e0b65";
		wait for Clk_period;
		Addr <=  "0001010001001";
		Trees_din <= x"5fff4604";
		wait for Clk_period;
		Addr <=  "0001010001010";
		Trees_din <= x"01f50b65";
		wait for Clk_period;
		Addr <=  "0001010001011";
		Trees_din <= x"00680b65";
		wait for Clk_period;
		Addr <=  "0001010001100";
		Trees_din <= x"ff830b65";
		wait for Clk_period;
		Addr <=  "0001010001101";
		Trees_din <= x"eaff4720";
		wait for Clk_period;
		Addr <=  "0001010001110";
		Trees_din <= x"76ffe710";
		wait for Clk_period;
		Addr <=  "0001010001111";
		Trees_din <= x"76ff6008";
		wait for Clk_period;
		Addr <=  "0001010010000";
		Trees_din <= x"4aff4904";
		wait for Clk_period;
		Addr <=  "0001010010001";
		Trees_din <= x"ffd10b65";
		wait for Clk_period;
		Addr <=  "0001010010010";
		Trees_din <= x"01630b65";
		wait for Clk_period;
		Addr <=  "0001010010011";
		Trees_din <= x"1afe5304";
		wait for Clk_period;
		Addr <=  "0001010010100";
		Trees_din <= x"00300b65";
		wait for Clk_period;
		Addr <=  "0001010010101";
		Trees_din <= x"ff630b65";
		wait for Clk_period;
		Addr <=  "0001010010110";
		Trees_din <= x"51007908";
		wait for Clk_period;
		Addr <=  "0001010010111";
		Trees_din <= x"a9fed804";
		wait for Clk_period;
		Addr <=  "0001010011000";
		Trees_din <= x"00da0b65";
		wait for Clk_period;
		Addr <=  "0001010011001";
		Trees_din <= x"ff9f0b65";
		wait for Clk_period;
		Addr <=  "0001010011010";
		Trees_din <= x"afff0604";
		wait for Clk_period;
		Addr <=  "0001010011011";
		Trees_din <= x"ffa40b65";
		wait for Clk_period;
		Addr <=  "0001010011100";
		Trees_din <= x"01640b65";
		wait for Clk_period;
		Addr <=  "0001010011101";
		Trees_din <= x"9dff4410";
		wait for Clk_period;
		Addr <=  "0001010011110";
		Trees_din <= x"c4002008";
		wait for Clk_period;
		Addr <=  "0001010011111";
		Trees_din <= x"73ff2404";
		wait for Clk_period;
		Addr <=  "0001010100000";
		Trees_din <= x"00aa0b65";
		wait for Clk_period;
		Addr <=  "0001010100001";
		Trees_din <= x"ff7b0b65";
		wait for Clk_period;
		Addr <=  "0001010100010";
		Trees_din <= x"87ff9604";
		wait for Clk_period;
		Addr <=  "0001010100011";
		Trees_din <= x"ffee0b65";
		wait for Clk_period;
		Addr <=  "0001010100100";
		Trees_din <= x"01300b65";
		wait for Clk_period;
		Addr <=  "0001010100101";
		Trees_din <= x"8effb508";
		wait for Clk_period;
		Addr <=  "0001010100110";
		Trees_din <= x"cb002f04";
		wait for Clk_period;
		Addr <=  "0001010100111";
		Trees_din <= x"00df0b65";
		wait for Clk_period;
		Addr <=  "0001010101000";
		Trees_din <= x"ffcc0b65";
		wait for Clk_period;
		Addr <=  "0001010101001";
		Trees_din <= x"91ffaa04";
		wait for Clk_period;
		Addr <=  "0001010101010";
		Trees_din <= x"005d0b65";
		wait for Clk_period;
		Addr <=  "0001010101011";
		Trees_din <= x"ffd50b65";
		wait for Clk_period;
		Addr <=  "0001010101100";
		Trees_din <= x"02fea72c";
		wait for Clk_period;
		Addr <=  "0001010101101";
		Trees_din <= x"5fff6f10";
		wait for Clk_period;
		Addr <=  "0001010101110";
		Trees_din <= x"a8ffbd0c";
		wait for Clk_period;
		Addr <=  "0001010101111";
		Trees_din <= x"5a00d208";
		wait for Clk_period;
		Addr <=  "0001010110000";
		Trees_din <= x"a4ffd704";
		wait for Clk_period;
		Addr <=  "0001010110001";
		Trees_din <= x"00d90b65";
		wait for Clk_period;
		Addr <=  "0001010110010";
		Trees_din <= x"ffdc0b65";
		wait for Clk_period;
		Addr <=  "0001010110011";
		Trees_din <= x"ff7e0b65";
		wait for Clk_period;
		Addr <=  "0001010110100";
		Trees_din <= x"ff710b65";
		wait for Clk_period;
		Addr <=  "0001010110101";
		Trees_din <= x"77fefe0c";
		wait for Clk_period;
		Addr <=  "0001010110110";
		Trees_din <= x"84ffe004";
		wait for Clk_period;
		Addr <=  "0001010110111";
		Trees_din <= x"ff820b65";
		wait for Clk_period;
		Addr <=  "0001010111000";
		Trees_din <= x"e5fe3304";
		wait for Clk_period;
		Addr <=  "0001010111001";
		Trees_din <= x"fff20b65";
		wait for Clk_period;
		Addr <=  "0001010111010";
		Trees_din <= x"01420b65";
		wait for Clk_period;
		Addr <=  "0001010111011";
		Trees_din <= x"55ffed08";
		wait for Clk_period;
		Addr <=  "0001010111100";
		Trees_din <= x"0dff6304";
		wait for Clk_period;
		Addr <=  "0001010111101";
		Trees_din <= x"00840b65";
		wait for Clk_period;
		Addr <=  "0001010111110";
		Trees_din <= x"00000b65";
		wait for Clk_period;
		Addr <=  "0001010111111";
		Trees_din <= x"3cfeb104";
		wait for Clk_period;
		Addr <=  "0001011000000";
		Trees_din <= x"00590b65";
		wait for Clk_period;
		Addr <=  "0001011000001";
		Trees_din <= x"02290b65";
		wait for Clk_period;
		Addr <=  "0001011000010";
		Trees_din <= x"56ff5b1c";
		wait for Clk_period;
		Addr <=  "0001011000011";
		Trees_din <= x"8e004610";
		wait for Clk_period;
		Addr <=  "0001011000100";
		Trees_din <= x"93ffbc08";
		wait for Clk_period;
		Addr <=  "0001011000101";
		Trees_din <= x"db007204";
		wait for Clk_period;
		Addr <=  "0001011000110";
		Trees_din <= x"ff8e0b65";
		wait for Clk_period;
		Addr <=  "0001011000111";
		Trees_din <= x"006f0b65";
		wait for Clk_period;
		Addr <=  "0001011001000";
		Trees_din <= x"9cff4504";
		wait for Clk_period;
		Addr <=  "0001011001001";
		Trees_din <= x"ff940b65";
		wait for Clk_period;
		Addr <=  "0001011001010";
		Trees_din <= x"00e50b65";
		wait for Clk_period;
		Addr <=  "0001011001011";
		Trees_din <= x"03011c08";
		wait for Clk_period;
		Addr <=  "0001011001100";
		Trees_din <= x"13017704";
		wait for Clk_period;
		Addr <=  "0001011001101";
		Trees_din <= x"ff680b65";
		wait for Clk_period;
		Addr <=  "0001011001110";
		Trees_din <= x"fff50b65";
		wait for Clk_period;
		Addr <=  "0001011001111";
		Trees_din <= x"00780b65";
		wait for Clk_period;
		Addr <=  "0001011010000";
		Trees_din <= x"0700f708";
		wait for Clk_period;
		Addr <=  "0001011010001";
		Trees_din <= x"a3006504";
		wait for Clk_period;
		Addr <=  "0001011010010";
		Trees_din <= x"ff5d0b65";
		wait for Clk_period;
		Addr <=  "0001011010011";
		Trees_din <= x"00570b65";
		wait for Clk_period;
		Addr <=  "0001011010100";
		Trees_din <= x"d5ffe704";
		wait for Clk_period;
		Addr <=  "0001011010101";
		Trees_din <= x"ff9b0b65";
		wait for Clk_period;
		Addr <=  "0001011010110";
		Trees_din <= x"0efe7504";
		wait for Clk_period;
		Addr <=  "0001011010111";
		Trees_din <= x"005a0b65";
		wait for Clk_period;
		Addr <=  "0001011011000";
		Trees_din <= x"01250b65";
		wait for Clk_period;
		Addr <=  "0001011011001";
		Trees_din <= x"19ffa078";
		wait for Clk_period;
		Addr <=  "0001011011010";
		Trees_din <= x"00ffa240";
		wait for Clk_period;
		Addr <=  "0001011011011";
		Trees_din <= x"4effef20";
		wait for Clk_period;
		Addr <=  "0001011011100";
		Trees_din <= x"76ffc910";
		wait for Clk_period;
		Addr <=  "0001011011101";
		Trees_din <= x"fefffc08";
		wait for Clk_period;
		Addr <=  "0001011011110";
		Trees_din <= x"20fff704";
		wait for Clk_period;
		Addr <=  "0001011011111";
		Trees_din <= x"ff9f0cd1";
		wait for Clk_period;
		Addr <=  "0001011100000";
		Trees_din <= x"000c0cd1";
		wait for Clk_period;
		Addr <=  "0001011100001";
		Trees_din <= x"2cffe304";
		wait for Clk_period;
		Addr <=  "0001011100010";
		Trees_din <= x"008b0cd1";
		wait for Clk_period;
		Addr <=  "0001011100011";
		Trees_din <= x"ffb30cd1";
		wait for Clk_period;
		Addr <=  "0001011100100";
		Trees_din <= x"8cffdb08";
		wait for Clk_period;
		Addr <=  "0001011100101";
		Trees_din <= x"41ff4404";
		wait for Clk_period;
		Addr <=  "0001011100110";
		Trees_din <= x"ffba0cd1";
		wait for Clk_period;
		Addr <=  "0001011100111";
		Trees_din <= x"004c0cd1";
		wait for Clk_period;
		Addr <=  "0001011101000";
		Trees_din <= x"b2ff8e04";
		wait for Clk_period;
		Addr <=  "0001011101001";
		Trees_din <= x"ffd40cd1";
		wait for Clk_period;
		Addr <=  "0001011101010";
		Trees_din <= x"007c0cd1";
		wait for Clk_period;
		Addr <=  "0001011101011";
		Trees_din <= x"04007410";
		wait for Clk_period;
		Addr <=  "0001011101100";
		Trees_din <= x"bbff7808";
		wait for Clk_period;
		Addr <=  "0001011101101";
		Trees_din <= x"03ff2704";
		wait for Clk_period;
		Addr <=  "0001011101110";
		Trees_din <= x"ff9b0cd1";
		wait for Clk_period;
		Addr <=  "0001011101111";
		Trees_din <= x"01130cd1";
		wait for Clk_period;
		Addr <=  "0001011110000";
		Trees_din <= x"01feac04";
		wait for Clk_period;
		Addr <=  "0001011110001";
		Trees_din <= x"00800cd1";
		wait for Clk_period;
		Addr <=  "0001011110010";
		Trees_din <= x"ff770cd1";
		wait for Clk_period;
		Addr <=  "0001011110011";
		Trees_din <= x"3dffd808";
		wait for Clk_period;
		Addr <=  "0001011110100";
		Trees_din <= x"85008204";
		wait for Clk_period;
		Addr <=  "0001011110101";
		Trees_din <= x"ff7b0cd1";
		wait for Clk_period;
		Addr <=  "0001011110110";
		Trees_din <= x"00780cd1";
		wait for Clk_period;
		Addr <=  "0001011110111";
		Trees_din <= x"d9ffdb04";
		wait for Clk_period;
		Addr <=  "0001011111000";
		Trees_din <= x"ffe50cd1";
		wait for Clk_period;
		Addr <=  "0001011111001";
		Trees_din <= x"00ef0cd1";
		wait for Clk_period;
		Addr <=  "0001011111010";
		Trees_din <= x"f4ff3818";
		wait for Clk_period;
		Addr <=  "0001011111011";
		Trees_din <= x"cd004810";
		wait for Clk_period;
		Addr <=  "0001011111100";
		Trees_din <= x"9a004008";
		wait for Clk_period;
		Addr <=  "0001011111101";
		Trees_din <= x"cf00c104";
		wait for Clk_period;
		Addr <=  "0001011111110";
		Trees_din <= x"008b0cd1";
		wait for Clk_period;
		Addr <=  "0001011111111";
		Trees_din <= x"ff720cd1";
		wait for Clk_period;
		Addr <=  "0001100000000";
		Trees_din <= x"8fff8004";
		wait for Clk_period;
		Addr <=  "0001100000001";
		Trees_din <= x"ff670cd1";
		wait for Clk_period;
		Addr <=  "0001100000010";
		Trees_din <= x"009d0cd1";
		wait for Clk_period;
		Addr <=  "0001100000011";
		Trees_din <= x"1f008004";
		wait for Clk_period;
		Addr <=  "0001100000100";
		Trees_din <= x"ff680cd1";
		wait for Clk_period;
		Addr <=  "0001100000101";
		Trees_din <= x"008b0cd1";
		wait for Clk_period;
		Addr <=  "0001100000110";
		Trees_din <= x"09000310";
		wait for Clk_period;
		Addr <=  "0001100000111";
		Trees_din <= x"93000208";
		wait for Clk_period;
		Addr <=  "0001100001000";
		Trees_din <= x"b9ffbc04";
		wait for Clk_period;
		Addr <=  "0001100001001";
		Trees_din <= x"ff7d0cd1";
		wait for Clk_period;
		Addr <=  "0001100001010";
		Trees_din <= x"007e0cd1";
		wait for Clk_period;
		Addr <=  "0001100001011";
		Trees_din <= x"fdff8504";
		wait for Clk_period;
		Addr <=  "0001100001100";
		Trees_din <= x"009c0cd1";
		wait for Clk_period;
		Addr <=  "0001100001101";
		Trees_din <= x"ff820cd1";
		wait for Clk_period;
		Addr <=  "0001100001110";
		Trees_din <= x"acffda08";
		wait for Clk_period;
		Addr <=  "0001100001111";
		Trees_din <= x"75009e04";
		wait for Clk_period;
		Addr <=  "0001100010000";
		Trees_din <= x"ff710cd1";
		wait for Clk_period;
		Addr <=  "0001100010001";
		Trees_din <= x"00560cd1";
		wait for Clk_period;
		Addr <=  "0001100010010";
		Trees_din <= x"88ff8b04";
		wait for Clk_period;
		Addr <=  "0001100010011";
		Trees_din <= x"ff9b0cd1";
		wait for Clk_period;
		Addr <=  "0001100010100";
		Trees_din <= x"00c90cd1";
		wait for Clk_period;
		Addr <=  "0001100010101";
		Trees_din <= x"db008d18";
		wait for Clk_period;
		Addr <=  "0001100010110";
		Trees_din <= x"dc007a0c";
		wait for Clk_period;
		Addr <=  "0001100010111";
		Trees_din <= x"4400ce08";
		wait for Clk_period;
		Addr <=  "0001100011000";
		Trees_din <= x"6bff7e04";
		wait for Clk_period;
		Addr <=  "0001100011001";
		Trees_din <= x"ff5b0cd1";
		wait for Clk_period;
		Addr <=  "0001100011010";
		Trees_din <= x"fff90cd1";
		wait for Clk_period;
		Addr <=  "0001100011011";
		Trees_din <= x"007e0cd1";
		wait for Clk_period;
		Addr <=  "0001100011100";
		Trees_din <= x"2bff5f08";
		wait for Clk_period;
		Addr <=  "0001100011101";
		Trees_din <= x"55001204";
		wait for Clk_period;
		Addr <=  "0001100011110";
		Trees_din <= x"01470cd1";
		wait for Clk_period;
		Addr <=  "0001100011111";
		Trees_din <= x"00020cd1";
		wait for Clk_period;
		Addr <=  "0001100100000";
		Trees_din <= x"ff7d0cd1";
		wait for Clk_period;
		Addr <=  "0001100100001";
		Trees_din <= x"b1fecc10";
		wait for Clk_period;
		Addr <=  "0001100100010";
		Trees_din <= x"16fea704";
		wait for Clk_period;
		Addr <=  "0001100100011";
		Trees_din <= x"ff8e0cd1";
		wait for Clk_period;
		Addr <=  "0001100100100";
		Trees_din <= x"7dffb604";
		wait for Clk_period;
		Addr <=  "0001100100101";
		Trees_din <= x"ffed0cd1";
		wait for Clk_period;
		Addr <=  "0001100100110";
		Trees_din <= x"5a009f04";
		wait for Clk_period;
		Addr <=  "0001100100111";
		Trees_din <= x"01980cd1";
		wait for Clk_period;
		Addr <=  "0001100101000";
		Trees_din <= x"002a0cd1";
		wait for Clk_period;
		Addr <=  "0001100101001";
		Trees_din <= x"34ffc308";
		wait for Clk_period;
		Addr <=  "0001100101010";
		Trees_din <= x"45ff2f04";
		wait for Clk_period;
		Addr <=  "0001100101011";
		Trees_din <= x"000d0cd1";
		wait for Clk_period;
		Addr <=  "0001100101100";
		Trees_din <= x"00ee0cd1";
		wait for Clk_period;
		Addr <=  "0001100101101";
		Trees_din <= x"16ff7308";
		wait for Clk_period;
		Addr <=  "0001100101110";
		Trees_din <= x"5100b604";
		wait for Clk_period;
		Addr <=  "0001100101111";
		Trees_din <= x"ff5f0cd1";
		wait for Clk_period;
		Addr <=  "0001100110000";
		Trees_din <= x"002f0cd1";
		wait for Clk_period;
		Addr <=  "0001100110001";
		Trees_din <= x"faffa204";
		wait for Clk_period;
		Addr <=  "0001100110010";
		Trees_din <= x"ffa30cd1";
		wait for Clk_period;
		Addr <=  "0001100110011";
		Trees_din <= x"00bc0cd1";
		wait for Clk_period;
		Addr <=  "0001100110100";
		Trees_din <= x"01fe7b64";
		wait for Clk_period;
		Addr <=  "0001100110101";
		Trees_din <= x"9bff723c";
		wait for Clk_period;
		Addr <=  "0001100110110";
		Trees_din <= x"e4fe561c";
		wait for Clk_period;
		Addr <=  "0001100110111";
		Trees_din <= x"6cffcf10";
		wait for Clk_period;
		Addr <=  "0001100111000";
		Trees_din <= x"51010608";
		wait for Clk_period;
		Addr <=  "0001100111001";
		Trees_din <= x"a2ff4b04";
		wait for Clk_period;
		Addr <=  "0001100111010";
		Trees_din <= x"004a0e0d";
		wait for Clk_period;
		Addr <=  "0001100111011";
		Trees_din <= x"ff900e0d";
		wait for Clk_period;
		Addr <=  "0001100111100";
		Trees_din <= x"d600d504";
		wait for Clk_period;
		Addr <=  "0001100111101";
		Trees_din <= x"ffe10e0d";
		wait for Clk_period;
		Addr <=  "0001100111110";
		Trees_din <= x"00b50e0d";
		wait for Clk_period;
		Addr <=  "0001100111111";
		Trees_din <= x"07009408";
		wait for Clk_period;
		Addr <=  "0001101000000";
		Trees_din <= x"8cff5e04";
		wait for Clk_period;
		Addr <=  "0001101000001";
		Trees_din <= x"ffd30e0d";
		wait for Clk_period;
		Addr <=  "0001101000010";
		Trees_din <= x"01010e0d";
		wait for Clk_period;
		Addr <=  "0001101000011";
		Trees_din <= x"ff7a0e0d";
		wait for Clk_period;
		Addr <=  "0001101000100";
		Trees_din <= x"71fedb10";
		wait for Clk_period;
		Addr <=  "0001101000101";
		Trees_din <= x"d9ffe608";
		wait for Clk_period;
		Addr <=  "0001101000110";
		Trees_din <= x"39fecb04";
		wait for Clk_period;
		Addr <=  "0001101000111";
		Trees_din <= x"00ae0e0d";
		wait for Clk_period;
		Addr <=  "0001101001000";
		Trees_din <= x"ffb00e0d";
		wait for Clk_period;
		Addr <=  "0001101001001";
		Trees_din <= x"2fff7904";
		wait for Clk_period;
		Addr <=  "0001101001010";
		Trees_din <= x"ffa30e0d";
		wait for Clk_period;
		Addr <=  "0001101001011";
		Trees_din <= x"00bd0e0d";
		wait for Clk_period;
		Addr <=  "0001101001100";
		Trees_din <= x"91000408";
		wait for Clk_period;
		Addr <=  "0001101001101";
		Trees_din <= x"7afef304";
		wait for Clk_period;
		Addr <=  "0001101001110";
		Trees_din <= x"ff7d0e0d";
		wait for Clk_period;
		Addr <=  "0001101001111";
		Trees_din <= x"00980e0d";
		wait for Clk_period;
		Addr <=  "0001101010000";
		Trees_din <= x"79ff0104";
		wait for Clk_period;
		Addr <=  "0001101010001";
		Trees_din <= x"000b0e0d";
		wait for Clk_period;
		Addr <=  "0001101010010";
		Trees_din <= x"ff730e0d";
		wait for Clk_period;
		Addr <=  "0001101010011";
		Trees_din <= x"56ffce20";
		wait for Clk_period;
		Addr <=  "0001101010100";
		Trees_din <= x"baffec10";
		wait for Clk_period;
		Addr <=  "0001101010101";
		Trees_din <= x"71fef808";
		wait for Clk_period;
		Addr <=  "0001101010110";
		Trees_din <= x"80ff3604";
		wait for Clk_period;
		Addr <=  "0001101010111";
		Trees_din <= x"ffa30e0d";
		wait for Clk_period;
		Addr <=  "0001101011000";
		Trees_din <= x"00c70e0d";
		wait for Clk_period;
		Addr <=  "0001101011001";
		Trees_din <= x"79fff604";
		wait for Clk_period;
		Addr <=  "0001101011010";
		Trees_din <= x"ffbb0e0d";
		wait for Clk_period;
		Addr <=  "0001101011011";
		Trees_din <= x"011a0e0d";
		wait for Clk_period;
		Addr <=  "0001101011100";
		Trees_din <= x"ebfe7208";
		wait for Clk_period;
		Addr <=  "0001101011101";
		Trees_din <= x"ceff8404";
		wait for Clk_period;
		Addr <=  "0001101011110";
		Trees_din <= x"011b0e0d";
		wait for Clk_period;
		Addr <=  "0001101011111";
		Trees_din <= x"ff920e0d";
		wait for Clk_period;
		Addr <=  "0001101100000";
		Trees_din <= x"db00f404";
		wait for Clk_period;
		Addr <=  "0001101100001";
		Trees_din <= x"ff610e0d";
		wait for Clk_period;
		Addr <=  "0001101100010";
		Trees_din <= x"00320e0d";
		wait for Clk_period;
		Addr <=  "0001101100011";
		Trees_din <= x"b4ff9504";
		wait for Clk_period;
		Addr <=  "0001101100100";
		Trees_din <= x"ff650e0d";
		wait for Clk_period;
		Addr <=  "0001101100101";
		Trees_din <= x"000f0e0d";
		wait for Clk_period;
		Addr <=  "0001101100110";
		Trees_din <= x"bbfff934";
		wait for Clk_period;
		Addr <=  "0001101100111";
		Trees_din <= x"19ffa020";
		wait for Clk_period;
		Addr <=  "0001101101000";
		Trees_din <= x"a4ff5810";
		wait for Clk_period;
		Addr <=  "0001101101001";
		Trees_din <= x"49ff6c08";
		wait for Clk_period;
		Addr <=  "0001101101010";
		Trees_din <= x"57ff2104";
		wait for Clk_period;
		Addr <=  "0001101101011";
		Trees_din <= x"01400e0d";
		wait for Clk_period;
		Addr <=  "0001101101100";
		Trees_din <= x"00200e0d";
		wait for Clk_period;
		Addr <=  "0001101101101";
		Trees_din <= x"a9febf04";
		wait for Clk_period;
		Addr <=  "0001101101110";
		Trees_din <= x"00fb0e0d";
		wait for Clk_period;
		Addr <=  "0001101101111";
		Trees_din <= x"000e0e0d";
		wait for Clk_period;
		Addr <=  "0001101110000";
		Trees_din <= x"5a00b608";
		wait for Clk_period;
		Addr <=  "0001101110001";
		Trees_din <= x"55001d04";
		wait for Clk_period;
		Addr <=  "0001101110010";
		Trees_din <= x"ffe00e0d";
		wait for Clk_period;
		Addr <=  "0001101110011";
		Trees_din <= x"003c0e0d";
		wait for Clk_period;
		Addr <=  "0001101110100";
		Trees_din <= x"b6ff8e04";
		wait for Clk_period;
		Addr <=  "0001101110101";
		Trees_din <= x"ff8e0e0d";
		wait for Clk_period;
		Addr <=  "0001101110110";
		Trees_din <= x"00120e0d";
		wait for Clk_period;
		Addr <=  "0001101110111";
		Trees_din <= x"ea004110";
		wait for Clk_period;
		Addr <=  "0001101111000";
		Trees_din <= x"79fed708";
		wait for Clk_period;
		Addr <=  "0001101111001";
		Trees_din <= x"f1ff5c04";
		wait for Clk_period;
		Addr <=  "0001101111010";
		Trees_din <= x"00d80e0d";
		wait for Clk_period;
		Addr <=  "0001101111011";
		Trees_din <= x"ffa10e0d";
		wait for Clk_period;
		Addr <=  "0001101111100";
		Trees_din <= x"69fe9504";
		wait for Clk_period;
		Addr <=  "0001101111101";
		Trees_din <= x"00190e0d";
		wait for Clk_period;
		Addr <=  "0001101111110";
		Trees_din <= x"ff600e0d";
		wait for Clk_period;
		Addr <=  "0001101111111";
		Trees_din <= x"00b70e0d";
		wait for Clk_period;
		Addr <=  "0001110000000";
		Trees_din <= x"7bfe4504";
		wait for Clk_period;
		Addr <=  "0001110000001";
		Trees_din <= x"00280e0d";
		wait for Clk_period;
		Addr <=  "0001110000010";
		Trees_din <= x"ff600e0d";
		wait for Clk_period;
		Addr <=  "0001110000011";
		Trees_din <= x"1aff3550";
		wait for Clk_period;
		Addr <=  "0001110000100";
		Trees_din <= x"bbfff934";
		wait for Clk_period;
		Addr <=  "0001110000101";
		Trees_din <= x"56002120";
		wait for Clk_period;
		Addr <=  "0001110000110";
		Trees_din <= x"19ff9e10";
		wait for Clk_period;
		Addr <=  "0001110000111";
		Trees_din <= x"a3fed208";
		wait for Clk_period;
		Addr <=  "0001110001000";
		Trees_din <= x"ab005f04";
		wait for Clk_period;
		Addr <=  "0001110001001";
		Trees_din <= x"ff650f29";
		wait for Clk_period;
		Addr <=  "0001110001010";
		Trees_din <= x"001a0f29";
		wait for Clk_period;
		Addr <=  "0001110001011";
		Trees_din <= x"31ff4704";
		wait for Clk_period;
		Addr <=  "0001110001100";
		Trees_din <= x"fff10f29";
		wait for Clk_period;
		Addr <=  "0001110001101";
		Trees_din <= x"00410f29";
		wait for Clk_period;
		Addr <=  "0001110001110";
		Trees_din <= x"db008d08";
		wait for Clk_period;
		Addr <=  "0001110001111";
		Trees_din <= x"ea004104";
		wait for Clk_period;
		Addr <=  "0001110010000";
		Trees_din <= x"ff810f29";
		wait for Clk_period;
		Addr <=  "0001110010001";
		Trees_din <= x"00af0f29";
		wait for Clk_period;
		Addr <=  "0001110010010";
		Trees_din <= x"b1fec604";
		wait for Clk_period;
		Addr <=  "0001110010011";
		Trees_din <= x"00b40f29";
		wait for Clk_period;
		Addr <=  "0001110010100";
		Trees_din <= x"ffdf0f29";
		wait for Clk_period;
		Addr <=  "0001110010101";
		Trees_din <= x"c9ff2d04";
		wait for Clk_period;
		Addr <=  "0001110010110";
		Trees_din <= x"012c0f29";
		wait for Clk_period;
		Addr <=  "0001110010111";
		Trees_din <= x"69fea708";
		wait for Clk_period;
		Addr <=  "0001110011000";
		Trees_din <= x"b0ffa404";
		wait for Clk_period;
		Addr <=  "0001110011001";
		Trees_din <= x"ffa00f29";
		wait for Clk_period;
		Addr <=  "0001110011010";
		Trees_din <= x"01040f29";
		wait for Clk_period;
		Addr <=  "0001110011011";
		Trees_din <= x"91fed204";
		wait for Clk_period;
		Addr <=  "0001110011100";
		Trees_din <= x"00710f29";
		wait for Clk_period;
		Addr <=  "0001110011101";
		Trees_din <= x"ff700f29";
		wait for Clk_period;
		Addr <=  "0001110011110";
		Trees_din <= x"a1002618";
		wait for Clk_period;
		Addr <=  "0001110011111";
		Trees_din <= x"31011110";
		wait for Clk_period;
		Addr <=  "0001110100000";
		Trees_din <= x"4dfdd408";
		wait for Clk_period;
		Addr <=  "0001110100001";
		Trees_din <= x"22ff4c04";
		wait for Clk_period;
		Addr <=  "0001110100010";
		Trees_din <= x"009f0f29";
		wait for Clk_period;
		Addr <=  "0001110100011";
		Trees_din <= x"ff9b0f29";
		wait for Clk_period;
		Addr <=  "0001110100100";
		Trees_din <= x"2b00da04";
		wait for Clk_period;
		Addr <=  "0001110100101";
		Trees_din <= x"ff5f0f29";
		wait for Clk_period;
		Addr <=  "0001110100110";
		Trees_din <= x"00050f29";
		wait for Clk_period;
		Addr <=  "0001110100111";
		Trees_din <= x"67ff2704";
		wait for Clk_period;
		Addr <=  "0001110101000";
		Trees_din <= x"ff9f0f29";
		wait for Clk_period;
		Addr <=  "0001110101001";
		Trees_din <= x"009b0f29";
		wait for Clk_period;
		Addr <=  "0001110101010";
		Trees_din <= x"00ba0f29";
		wait for Clk_period;
		Addr <=  "0001110101011";
		Trees_din <= x"1bff7910";
		wait for Clk_period;
		Addr <=  "0001110101100";
		Trees_din <= x"8800ae08";
		wait for Clk_period;
		Addr <=  "0001110101101";
		Trees_din <= x"7f002504";
		wait for Clk_period;
		Addr <=  "0001110101110";
		Trees_din <= x"ff610f29";
		wait for Clk_period;
		Addr <=  "0001110101111";
		Trees_din <= x"00360f29";
		wait for Clk_period;
		Addr <=  "0001110110000";
		Trees_din <= x"25002904";
		wait for Clk_period;
		Addr <=  "0001110110001";
		Trees_din <= x"00160f29";
		wait for Clk_period;
		Addr <=  "0001110110010";
		Trees_din <= x"00a90f29";
		wait for Clk_period;
		Addr <=  "0001110110011";
		Trees_din <= x"a5feb014";
		wait for Clk_period;
		Addr <=  "0001110110100";
		Trees_din <= x"dcff9d04";
		wait for Clk_period;
		Addr <=  "0001110110101";
		Trees_din <= x"ff860f29";
		wait for Clk_period;
		Addr <=  "0001110110110";
		Trees_din <= x"90ffbe08";
		wait for Clk_period;
		Addr <=  "0001110110111";
		Trees_din <= x"c2ff8704";
		wait for Clk_period;
		Addr <=  "0001110111000";
		Trees_din <= x"018d0f29";
		wait for Clk_period;
		Addr <=  "0001110111001";
		Trees_din <= x"00050f29";
		wait for Clk_period;
		Addr <=  "0001110111010";
		Trees_din <= x"eaffa704";
		wait for Clk_period;
		Addr <=  "0001110111011";
		Trees_din <= x"ffac0f29";
		wait for Clk_period;
		Addr <=  "0001110111100";
		Trees_din <= x"00110f29";
		wait for Clk_period;
		Addr <=  "0001110111101";
		Trees_din <= x"9efed40c";
		wait for Clk_period;
		Addr <=  "0001110111110";
		Trees_din <= x"b1fee704";
		wait for Clk_period;
		Addr <=  "0001110111111";
		Trees_din <= x"01880f29";
		wait for Clk_period;
		Addr <=  "0001111000000";
		Trees_din <= x"6e00ca04";
		wait for Clk_period;
		Addr <=  "0001111000001";
		Trees_din <= x"ff910f29";
		wait for Clk_period;
		Addr <=  "0001111000010";
		Trees_din <= x"00a40f29";
		wait for Clk_period;
		Addr <=  "0001111000011";
		Trees_din <= x"39ffa008";
		wait for Clk_period;
		Addr <=  "0001111000100";
		Trees_din <= x"57fec304";
		wait for Clk_period;
		Addr <=  "0001111000101";
		Trees_din <= x"009c0f29";
		wait for Clk_period;
		Addr <=  "0001111000110";
		Trees_din <= x"ffcf0f29";
		wait for Clk_period;
		Addr <=  "0001111000111";
		Trees_din <= x"a9fec304";
		wait for Clk_period;
		Addr <=  "0001111001000";
		Trees_din <= x"00b40f29";
		wait for Clk_period;
		Addr <=  "0001111001001";
		Trees_din <= x"ff830f29";
		wait for Clk_period;
		Addr <=  "0001111001010";
		Trees_din <= x"fcfebd38";
		wait for Clk_period;
		Addr <=  "0001111001011";
		Trees_din <= x"1fffba0c";
		wait for Clk_period;
		Addr <=  "0001111001100";
		Trees_din <= x"0b006304";
		wait for Clk_period;
		Addr <=  "0001111001101";
		Trees_din <= x"ff601085";
		wait for Clk_period;
		Addr <=  "0001111001110";
		Trees_din <= x"40ffeb04";
		wait for Clk_period;
		Addr <=  "0001111001111";
		Trees_din <= x"00961085";
		wait for Clk_period;
		Addr <=  "0001111010000";
		Trees_din <= x"ff871085";
		wait for Clk_period;
		Addr <=  "0001111010001";
		Trees_din <= x"fdffb518";
		wait for Clk_period;
		Addr <=  "0001111010010";
		Trees_din <= x"35fe330c";
		wait for Clk_period;
		Addr <=  "0001111010011";
		Trees_din <= x"36ff7108";
		wait for Clk_period;
		Addr <=  "0001111010100";
		Trees_din <= x"deffff04";
		wait for Clk_period;
		Addr <=  "0001111010101";
		Trees_din <= x"ffa61085";
		wait for Clk_period;
		Addr <=  "0001111010110";
		Trees_din <= x"00091085";
		wait for Clk_period;
		Addr <=  "0001111010111";
		Trees_din <= x"00cd1085";
		wait for Clk_period;
		Addr <=  "0001111011000";
		Trees_din <= x"00002408";
		wait for Clk_period;
		Addr <=  "0001111011001";
		Trees_din <= x"aaff2004";
		wait for Clk_period;
		Addr <=  "0001111011010";
		Trees_din <= x"00081085";
		wait for Clk_period;
		Addr <=  "0001111011011";
		Trees_din <= x"ff651085";
		wait for Clk_period;
		Addr <=  "0001111011100";
		Trees_din <= x"00841085";
		wait for Clk_period;
		Addr <=  "0001111011101";
		Trees_din <= x"7dff8e04";
		wait for Clk_period;
		Addr <=  "0001111011110";
		Trees_din <= x"ff861085";
		wait for Clk_period;
		Addr <=  "0001111011111";
		Trees_din <= x"9eff1c08";
		wait for Clk_period;
		Addr <=  "0001111100000";
		Trees_din <= x"65ff0d04";
		wait for Clk_period;
		Addr <=  "0001111100001";
		Trees_din <= x"ffa01085";
		wait for Clk_period;
		Addr <=  "0001111100010";
		Trees_din <= x"fff41085";
		wait for Clk_period;
		Addr <=  "0001111100011";
		Trees_din <= x"87ff3a04";
		wait for Clk_period;
		Addr <=  "0001111100100";
		Trees_din <= x"00151085";
		wait for Clk_period;
		Addr <=  "0001111100101";
		Trees_din <= x"012d1085";
		wait for Clk_period;
		Addr <=  "0001111100110";
		Trees_din <= x"b1ff1440";
		wait for Clk_period;
		Addr <=  "0001111100111";
		Trees_din <= x"36ffcb20";
		wait for Clk_period;
		Addr <=  "0001111101000";
		Trees_din <= x"c9ffb710";
		wait for Clk_period;
		Addr <=  "0001111101001";
		Trees_din <= x"6c005608";
		wait for Clk_period;
		Addr <=  "0001111101010";
		Trees_din <= x"e9ff0b04";
		wait for Clk_period;
		Addr <=  "0001111101011";
		Trees_din <= x"001f1085";
		wait for Clk_period;
		Addr <=  "0001111101100";
		Trees_din <= x"ffb01085";
		wait for Clk_period;
		Addr <=  "0001111101101";
		Trees_din <= x"21ff8904";
		wait for Clk_period;
		Addr <=  "0001111101110";
		Trees_din <= x"01701085";
		wait for Clk_period;
		Addr <=  "0001111101111";
		Trees_din <= x"fff81085";
		wait for Clk_period;
		Addr <=  "0001111110000";
		Trees_din <= x"90ff4508";
		wait for Clk_period;
		Addr <=  "0001111110001";
		Trees_din <= x"89008204";
		wait for Clk_period;
		Addr <=  "0001111110010";
		Trees_din <= x"fff51085";
		wait for Clk_period;
		Addr <=  "0001111110011";
		Trees_din <= x"009a1085";
		wait for Clk_period;
		Addr <=  "0001111110100";
		Trees_din <= x"b3fe8404";
		wait for Clk_period;
		Addr <=  "0001111110101";
		Trees_din <= x"ffa31085";
		wait for Clk_period;
		Addr <=  "0001111110110";
		Trees_din <= x"00861085";
		wait for Clk_period;
		Addr <=  "0001111110111";
		Trees_din <= x"20005a10";
		wait for Clk_period;
		Addr <=  "0001111111000";
		Trees_din <= x"be007b08";
		wait for Clk_period;
		Addr <=  "0001111111001";
		Trees_din <= x"4effd704";
		wait for Clk_period;
		Addr <=  "0001111111010";
		Trees_din <= x"ff701085";
		wait for Clk_period;
		Addr <=  "0001111111011";
		Trees_din <= x"00241085";
		wait for Clk_period;
		Addr <=  "0001111111100";
		Trees_din <= x"5fff6604";
		wait for Clk_period;
		Addr <=  "0001111111101";
		Trees_din <= x"ff9b1085";
		wait for Clk_period;
		Addr <=  "0001111111110";
		Trees_din <= x"00e71085";
		wait for Clk_period;
		Addr <=  "0001111111111";
		Trees_din <= x"c2ff8b08";
		wait for Clk_period;
		Addr <=  "0010000000000";
		Trees_din <= x"c8006804";
		wait for Clk_period;
		Addr <=  "0010000000001";
		Trees_din <= x"ff991085";
		wait for Clk_period;
		Addr <=  "0010000000010";
		Trees_din <= x"00391085";
		wait for Clk_period;
		Addr <=  "0010000000011";
		Trees_din <= x"aaff7704";
		wait for Clk_period;
		Addr <=  "0010000000100";
		Trees_din <= x"00331085";
		wait for Clk_period;
		Addr <=  "0010000000101";
		Trees_din <= x"00e21085";
		wait for Clk_period;
		Addr <=  "0010000000110";
		Trees_din <= x"6d00241c";
		wait for Clk_period;
		Addr <=  "0010000000111";
		Trees_din <= x"e6000310";
		wait for Clk_period;
		Addr <=  "0010000001000";
		Trees_din <= x"36ff7c08";
		wait for Clk_period;
		Addr <=  "0010000001001";
		Trees_din <= x"56ff8b04";
		wait for Clk_period;
		Addr <=  "0010000001010";
		Trees_din <= x"002c1085";
		wait for Clk_period;
		Addr <=  "0010000001011";
		Trees_din <= x"ffb51085";
		wait for Clk_period;
		Addr <=  "0010000001100";
		Trees_din <= x"2efeac04";
		wait for Clk_period;
		Addr <=  "0010000001101";
		Trees_din <= x"009a1085";
		wait for Clk_period;
		Addr <=  "0010000001110";
		Trees_din <= x"ff891085";
		wait for Clk_period;
		Addr <=  "0010000001111";
		Trees_din <= x"8e00dd08";
		wait for Clk_period;
		Addr <=  "0010000010000";
		Trees_din <= x"b5ff7f04";
		wait for Clk_period;
		Addr <=  "0010000010001";
		Trees_din <= x"ff5f1085";
		wait for Clk_period;
		Addr <=  "0010000010010";
		Trees_din <= x"fff31085";
		wait for Clk_period;
		Addr <=  "0010000010011";
		Trees_din <= x"00931085";
		wait for Clk_period;
		Addr <=  "0010000010100";
		Trees_din <= x"9dffe110";
		wait for Clk_period;
		Addr <=  "0010000010101";
		Trees_din <= x"f4fe6508";
		wait for Clk_period;
		Addr <=  "0010000010110";
		Trees_din <= x"9a000804";
		wait for Clk_period;
		Addr <=  "0010000010111";
		Trees_din <= x"00b71085";
		wait for Clk_period;
		Addr <=  "0010000011000";
		Trees_din <= x"ff7f1085";
		wait for Clk_period;
		Addr <=  "0010000011001";
		Trees_din <= x"2b004204";
		wait for Clk_period;
		Addr <=  "0010000011010";
		Trees_din <= x"ffd41085";
		wait for Clk_period;
		Addr <=  "0010000011011";
		Trees_din <= x"004b1085";
		wait for Clk_period;
		Addr <=  "0010000011100";
		Trees_din <= x"e4fe0604";
		wait for Clk_period;
		Addr <=  "0010000011101";
		Trees_din <= x"ff7d1085";
		wait for Clk_period;
		Addr <=  "0010000011110";
		Trees_din <= x"4afed104";
		wait for Clk_period;
		Addr <=  "0010000011111";
		Trees_din <= x"01121085";
		wait for Clk_period;
		Addr <=  "0010000100000";
		Trees_din <= x"004a1085";
		wait for Clk_period;
		Addr <=  "0010000100001";
		Trees_din <= x"01fe7f7c";
		wait for Clk_period;
		Addr <=  "0010000100010";
		Trees_din <= x"83ff3b3c";
		wait for Clk_period;
		Addr <=  "0010000100011";
		Trees_din <= x"b4feee1c";
		wait for Clk_period;
		Addr <=  "0010000100100";
		Trees_din <= x"1fff480c";
		wait for Clk_period;
		Addr <=  "0010000100101";
		Trees_din <= x"9eff0708";
		wait for Clk_period;
		Addr <=  "0010000100110";
		Trees_din <= x"feff4204";
		wait for Clk_period;
		Addr <=  "0010000100111";
		Trees_din <= x"00d21259";
		wait for Clk_period;
		Addr <=  "0010000101000";
		Trees_din <= x"ffae1259";
		wait for Clk_period;
		Addr <=  "0010000101001";
		Trees_din <= x"ff6c1259";
		wait for Clk_period;
		Addr <=  "0010000101010";
		Trees_din <= x"a4ffd808";
		wait for Clk_period;
		Addr <=  "0010000101011";
		Trees_din <= x"67ff4f04";
		wait for Clk_period;
		Addr <=  "0010000101100";
		Trees_din <= x"00821259";
		wait for Clk_period;
		Addr <=  "0010000101101";
		Trees_din <= x"00131259";
		wait for Clk_period;
		Addr <=  "0010000101110";
		Trees_din <= x"2aff9b04";
		wait for Clk_period;
		Addr <=  "0010000101111";
		Trees_din <= x"00021259";
		wait for Clk_period;
		Addr <=  "0010000110000";
		Trees_din <= x"ff761259";
		wait for Clk_period;
		Addr <=  "0010000110001";
		Trees_din <= x"ab00ac10";
		wait for Clk_period;
		Addr <=  "0010000110010";
		Trees_din <= x"e4fef008";
		wait for Clk_period;
		Addr <=  "0010000110011";
		Trees_din <= x"22fee504";
		wait for Clk_period;
		Addr <=  "0010000110100";
		Trees_din <= x"002d1259";
		wait for Clk_period;
		Addr <=  "0010000110101";
		Trees_din <= x"ff611259";
		wait for Clk_period;
		Addr <=  "0010000110110";
		Trees_din <= x"8aff5204";
		wait for Clk_period;
		Addr <=  "0010000110111";
		Trees_din <= x"00ec1259";
		wait for Clk_period;
		Addr <=  "0010000111000";
		Trees_din <= x"ffad1259";
		wait for Clk_period;
		Addr <=  "0010000111001";
		Trees_din <= x"d7005e08";
		wait for Clk_period;
		Addr <=  "0010000111010";
		Trees_din <= x"6bff4804";
		wait for Clk_period;
		Addr <=  "0010000111011";
		Trees_din <= x"ff751259";
		wait for Clk_period;
		Addr <=  "0010000111100";
		Trees_din <= x"003d1259";
		wait for Clk_period;
		Addr <=  "0010000111101";
		Trees_din <= x"c5ff3e04";
		wait for Clk_period;
		Addr <=  "0010000111110";
		Trees_din <= x"00a61259";
		wait for Clk_period;
		Addr <=  "0010000111111";
		Trees_din <= x"ffd71259";
		wait for Clk_period;
		Addr <=  "0010001000000";
		Trees_din <= x"25002420";
		wait for Clk_period;
		Addr <=  "0010001000001";
		Trees_din <= x"60ffba10";
		wait for Clk_period;
		Addr <=  "0010001000010";
		Trees_din <= x"16ff7808";
		wait for Clk_period;
		Addr <=  "0010001000011";
		Trees_din <= x"35fe7b04";
		wait for Clk_period;
		Addr <=  "0010001000100";
		Trees_din <= x"00151259";
		wait for Clk_period;
		Addr <=  "0010001000101";
		Trees_din <= x"00d01259";
		wait for Clk_period;
		Addr <=  "0010001000110";
		Trees_din <= x"0eff1104";
		wait for Clk_period;
		Addr <=  "0010001000111";
		Trees_din <= x"ff861259";
		wait for Clk_period;
		Addr <=  "0010001001000";
		Trees_din <= x"fffa1259";
		wait for Clk_period;
		Addr <=  "0010001001001";
		Trees_din <= x"e4fed808";
		wait for Clk_period;
		Addr <=  "0010001001010";
		Trees_din <= x"ceffdc04";
		wait for Clk_period;
		Addr <=  "0010001001011";
		Trees_din <= x"00d71259";
		wait for Clk_period;
		Addr <=  "0010001001100";
		Trees_din <= x"ffc21259";
		wait for Clk_period;
		Addr <=  "0010001001101";
		Trees_din <= x"5dffbc04";
		wait for Clk_period;
		Addr <=  "0010001001110";
		Trees_din <= x"ff6b1259";
		wait for Clk_period;
		Addr <=  "0010001001111";
		Trees_din <= x"ffeb1259";
		wait for Clk_period;
		Addr <=  "0010001010000";
		Trees_din <= x"9bff7010";
		wait for Clk_period;
		Addr <=  "0010001010001";
		Trees_din <= x"e1ffa408";
		wait for Clk_period;
		Addr <=  "0010001010010";
		Trees_din <= x"90ffbb04";
		wait for Clk_period;
		Addr <=  "0010001010011";
		Trees_din <= x"00c31259";
		wait for Clk_period;
		Addr <=  "0010001010100";
		Trees_din <= x"ff931259";
		wait for Clk_period;
		Addr <=  "0010001010101";
		Trees_din <= x"f1ff5304";
		wait for Clk_period;
		Addr <=  "0010001010110";
		Trees_din <= x"ff811259";
		wait for Clk_period;
		Addr <=  "0010001010111";
		Trees_din <= x"00391259";
		wait for Clk_period;
		Addr <=  "0010001011000";
		Trees_din <= x"68ff2e08";
		wait for Clk_period;
		Addr <=  "0010001011001";
		Trees_din <= x"d2fe5104";
		wait for Clk_period;
		Addr <=  "0010001011010";
		Trees_din <= x"00211259";
		wait for Clk_period;
		Addr <=  "0010001011011";
		Trees_din <= x"ff651259";
		wait for Clk_period;
		Addr <=  "0010001011100";
		Trees_din <= x"cdffa904";
		wait for Clk_period;
		Addr <=  "0010001011101";
		Trees_din <= x"00801259";
		wait for Clk_period;
		Addr <=  "0010001011110";
		Trees_din <= x"ffa81259";
		wait for Clk_period;
		Addr <=  "0010001011111";
		Trees_din <= x"6bfe9b30";
		wait for Clk_period;
		Addr <=  "0010001100000";
		Trees_din <= x"a9ffb620";
		wait for Clk_period;
		Addr <=  "0010001100001";
		Trees_din <= x"99ff1910";
		wait for Clk_period;
		Addr <=  "0010001100010";
		Trees_din <= x"bcffdc08";
		wait for Clk_period;
		Addr <=  "0010001100011";
		Trees_din <= x"02fea404";
		wait for Clk_period;
		Addr <=  "0010001100100";
		Trees_din <= x"ffe81259";
		wait for Clk_period;
		Addr <=  "0010001100101";
		Trees_din <= x"ff741259";
		wait for Clk_period;
		Addr <=  "0010001100110";
		Trees_din <= x"7aff6e04";
		wait for Clk_period;
		Addr <=  "0010001100111";
		Trees_din <= x"01171259";
		wait for Clk_period;
		Addr <=  "0010001101000";
		Trees_din <= x"001a1259";
		wait for Clk_period;
		Addr <=  "0010001101001";
		Trees_din <= x"6fff2e08";
		wait for Clk_period;
		Addr <=  "0010001101010";
		Trees_din <= x"faff6a04";
		wait for Clk_period;
		Addr <=  "0010001101011";
		Trees_din <= x"015d1259";
		wait for Clk_period;
		Addr <=  "0010001101100";
		Trees_din <= x"ffd91259";
		wait for Clk_period;
		Addr <=  "0010001101101";
		Trees_din <= x"d9ffaa04";
		wait for Clk_period;
		Addr <=  "0010001101110";
		Trees_din <= x"00671259";
		wait for Clk_period;
		Addr <=  "0010001101111";
		Trees_din <= x"ff9f1259";
		wait for Clk_period;
		Addr <=  "0010001110000";
		Trees_din <= x"8100480c";
		wait for Clk_period;
		Addr <=  "0010001110001";
		Trees_din <= x"e7004a08";
		wait for Clk_period;
		Addr <=  "0010001110010";
		Trees_din <= x"6ffeb704";
		wait for Clk_period;
		Addr <=  "0010001110011";
		Trees_din <= x"00191259";
		wait for Clk_period;
		Addr <=  "0010001110100";
		Trees_din <= x"ff601259";
		wait for Clk_period;
		Addr <=  "0010001110101";
		Trees_din <= x"00251259";
		wait for Clk_period;
		Addr <=  "0010001110110";
		Trees_din <= x"00351259";
		wait for Clk_period;
		Addr <=  "0010001110111";
		Trees_din <= x"10ffdb20";
		wait for Clk_period;
		Addr <=  "0010001111000";
		Trees_din <= x"37ffea10";
		wait for Clk_period;
		Addr <=  "0010001111001";
		Trees_din <= x"ac00a408";
		wait for Clk_period;
		Addr <=  "0010001111010";
		Trees_din <= x"b6ff7204";
		wait for Clk_period;
		Addr <=  "0010001111011";
		Trees_din <= x"ffc71259";
		wait for Clk_period;
		Addr <=  "0010001111100";
		Trees_din <= x"00241259";
		wait for Clk_period;
		Addr <=  "0010001111101";
		Trees_din <= x"0efe8904";
		wait for Clk_period;
		Addr <=  "0010001111110";
		Trees_din <= x"ffbc1259";
		wait for Clk_period;
		Addr <=  "0010001111111";
		Trees_din <= x"011c1259";
		wait for Clk_period;
		Addr <=  "0010010000000";
		Trees_din <= x"beff5c08";
		wait for Clk_period;
		Addr <=  "0010010000001";
		Trees_din <= x"1cff4104";
		wait for Clk_period;
		Addr <=  "0010010000010";
		Trees_din <= x"01331259";
		wait for Clk_period;
		Addr <=  "0010010000011";
		Trees_din <= x"ff9f1259";
		wait for Clk_period;
		Addr <=  "0010010000100";
		Trees_din <= x"61007a04";
		wait for Clk_period;
		Addr <=  "0010010000101";
		Trees_din <= x"ff661259";
		wait for Clk_period;
		Addr <=  "0010010000110";
		Trees_din <= x"00401259";
		wait for Clk_period;
		Addr <=  "0010010000111";
		Trees_din <= x"feff1310";
		wait for Clk_period;
		Addr <=  "0010010001000";
		Trees_din <= x"8ffeea08";
		wait for Clk_period;
		Addr <=  "0010010001001";
		Trees_din <= x"53ff8204";
		wait for Clk_period;
		Addr <=  "0010010001010";
		Trees_din <= x"01841259";
		wait for Clk_period;
		Addr <=  "0010010001011";
		Trees_din <= x"00791259";
		wait for Clk_period;
		Addr <=  "0010010001100";
		Trees_din <= x"51ffb804";
		wait for Clk_period;
		Addr <=  "0010010001101";
		Trees_din <= x"003c1259";
		wait for Clk_period;
		Addr <=  "0010010001110";
		Trees_din <= x"ffa71259";
		wait for Clk_period;
		Addr <=  "0010010001111";
		Trees_din <= x"feff9808";
		wait for Clk_period;
		Addr <=  "0010010010000";
		Trees_din <= x"4fffcc04";
		wait for Clk_period;
		Addr <=  "0010010010001";
		Trees_din <= x"ff8b1259";
		wait for Clk_period;
		Addr <=  "0010010010010";
		Trees_din <= x"00421259";
		wait for Clk_period;
		Addr <=  "0010010010011";
		Trees_din <= x"3cfebe04";
		wait for Clk_period;
		Addr <=  "0010010010100";
		Trees_din <= x"ffba1259";
		wait for Clk_period;
		Addr <=  "0010010010101";
		Trees_din <= x"00541259";
		wait for Clk_period;
		Addr <=  "0010010010110";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0010010010111";
		Trees_din <= x"19ffa058";
		wait for Clk_period;
		Addr <=  "0010010011000";
		Trees_din <= x"20feec20";
		wait for Clk_period;
		Addr <=  "0010010011001";
		Trees_din <= x"61007a1c";
		wait for Clk_period;
		Addr <=  "0010010011010";
		Trees_din <= x"b9ff940c";
		wait for Clk_period;
		Addr <=  "0010010011011";
		Trees_din <= x"93fff404";
		wait for Clk_period;
		Addr <=  "0010010011100";
		Trees_din <= x"ff631379";
		wait for Clk_period;
		Addr <=  "0010010011101";
		Trees_din <= x"5bff7f04";
		wait for Clk_period;
		Addr <=  "0010010011110";
		Trees_din <= x"ff8c1379";
		wait for Clk_period;
		Addr <=  "0010010011111";
		Trees_din <= x"00781379";
		wait for Clk_period;
		Addr <=  "0010010100000";
		Trees_din <= x"2aff8608";
		wait for Clk_period;
		Addr <=  "0010010100001";
		Trees_din <= x"1eff7104";
		wait for Clk_period;
		Addr <=  "0010010100010";
		Trees_din <= x"00f61379";
		wait for Clk_period;
		Addr <=  "0010010100011";
		Trees_din <= x"000a1379";
		wait for Clk_period;
		Addr <=  "0010010100100";
		Trees_din <= x"30000504";
		wait for Clk_period;
		Addr <=  "0010010100101";
		Trees_din <= x"ff911379";
		wait for Clk_period;
		Addr <=  "0010010100110";
		Trees_din <= x"fffa1379";
		wait for Clk_period;
		Addr <=  "0010010100111";
		Trees_din <= x"00c51379";
		wait for Clk_period;
		Addr <=  "0010010101000";
		Trees_din <= x"fcfebc18";
		wait for Clk_period;
		Addr <=  "0010010101001";
		Trees_din <= x"1fffba08";
		wait for Clk_period;
		Addr <=  "0010010101010";
		Trees_din <= x"2600d304";
		wait for Clk_period;
		Addr <=  "0010010101011";
		Trees_din <= x"ff641379";
		wait for Clk_period;
		Addr <=  "0010010101100";
		Trees_din <= x"00271379";
		wait for Clk_period;
		Addr <=  "0010010101101";
		Trees_din <= x"fdffb508";
		wait for Clk_period;
		Addr <=  "0010010101110";
		Trees_din <= x"d3fee104";
		wait for Clk_period;
		Addr <=  "0010010101111";
		Trees_din <= x"00181379";
		wait for Clk_period;
		Addr <=  "0010010110000";
		Trees_din <= x"ff7c1379";
		wait for Clk_period;
		Addr <=  "0010010110001";
		Trees_din <= x"9affad04";
		wait for Clk_period;
		Addr <=  "0010010110010";
		Trees_din <= x"00b31379";
		wait for Clk_period;
		Addr <=  "0010010110011";
		Trees_din <= x"ffd81379";
		wait for Clk_period;
		Addr <=  "0010010110100";
		Trees_din <= x"bbfff910";
		wait for Clk_period;
		Addr <=  "0010010110101";
		Trees_din <= x"b1ff1408";
		wait for Clk_period;
		Addr <=  "0010010110110";
		Trees_din <= x"89fef804";
		wait for Clk_period;
		Addr <=  "0010010110111";
		Trees_din <= x"ff6d1379";
		wait for Clk_period;
		Addr <=  "0010010111000";
		Trees_din <= x"00431379";
		wait for Clk_period;
		Addr <=  "0010010111001";
		Trees_din <= x"6d000904";
		wait for Clk_period;
		Addr <=  "0010010111010";
		Trees_din <= x"ffd81379";
		wait for Clk_period;
		Addr <=  "0010010111011";
		Trees_din <= x"00281379";
		wait for Clk_period;
		Addr <=  "0010010111100";
		Trees_din <= x"d2fe3308";
		wait for Clk_period;
		Addr <=  "0010010111101";
		Trees_din <= x"3bff3604";
		wait for Clk_period;
		Addr <=  "0010010111110";
		Trees_din <= x"00091379";
		wait for Clk_period;
		Addr <=  "0010010111111";
		Trees_din <= x"00951379";
		wait for Clk_period;
		Addr <=  "0010011000000";
		Trees_din <= x"4dfdd404";
		wait for Clk_period;
		Addr <=  "0010011000001";
		Trees_din <= x"00321379";
		wait for Clk_period;
		Addr <=  "0010011000010";
		Trees_din <= x"ff761379";
		wait for Clk_period;
		Addr <=  "0010011000011";
		Trees_din <= x"db008d18";
		wait for Clk_period;
		Addr <=  "0010011000100";
		Trees_din <= x"dc007a0c";
		wait for Clk_period;
		Addr <=  "0010011000101";
		Trees_din <= x"4400ce08";
		wait for Clk_period;
		Addr <=  "0010011000110";
		Trees_din <= x"30007e04";
		wait for Clk_period;
		Addr <=  "0010011000111";
		Trees_din <= x"ff621379";
		wait for Clk_period;
		Addr <=  "0010011001000";
		Trees_din <= x"fff81379";
		wait for Clk_period;
		Addr <=  "0010011001001";
		Trees_din <= x"004a1379";
		wait for Clk_period;
		Addr <=  "0010011001010";
		Trees_din <= x"2bff5f08";
		wait for Clk_period;
		Addr <=  "0010011001011";
		Trees_din <= x"6bfe8b04";
		wait for Clk_period;
		Addr <=  "0010011001100";
		Trees_din <= x"00081379";
		wait for Clk_period;
		Addr <=  "0010011001101";
		Trees_din <= x"00d91379";
		wait for Clk_period;
		Addr <=  "0010011001110";
		Trees_din <= x"ff8b1379";
		wait for Clk_period;
		Addr <=  "0010011001111";
		Trees_din <= x"e0fef308";
		wait for Clk_period;
		Addr <=  "0010011010000";
		Trees_din <= x"72007204";
		wait for Clk_period;
		Addr <=  "0010011010001";
		Trees_din <= x"ff731379";
		wait for Clk_period;
		Addr <=  "0010011010010";
		Trees_din <= x"003f1379";
		wait for Clk_period;
		Addr <=  "0010011010011";
		Trees_din <= x"3dffae08";
		wait for Clk_period;
		Addr <=  "0010011010100";
		Trees_din <= x"d4fee004";
		wait for Clk_period;
		Addr <=  "0010011010101";
		Trees_din <= x"00731379";
		wait for Clk_period;
		Addr <=  "0010011010110";
		Trees_din <= x"ff791379";
		wait for Clk_period;
		Addr <=  "0010011010111";
		Trees_din <= x"d5ffed08";
		wait for Clk_period;
		Addr <=  "0010011011000";
		Trees_din <= x"dfff9f04";
		wait for Clk_period;
		Addr <=  "0010011011001";
		Trees_din <= x"ff8f1379";
		wait for Clk_period;
		Addr <=  "0010011011010";
		Trees_din <= x"00761379";
		wait for Clk_period;
		Addr <=  "0010011011011";
		Trees_din <= x"a3ff3b04";
		wait for Clk_period;
		Addr <=  "0010011011100";
		Trees_din <= x"003f1379";
		wait for Clk_period;
		Addr <=  "0010011011101";
		Trees_din <= x"00f51379";
		wait for Clk_period;
		Addr <=  "0010011011110";
		Trees_din <= x"ab008e50";
		wait for Clk_period;
		Addr <=  "0010011011111";
		Trees_din <= x"7afef810";
		wait for Clk_period;
		Addr <=  "0010011100000";
		Trees_din <= x"b4fe4608";
		wait for Clk_period;
		Addr <=  "0010011100001";
		Trees_din <= x"10003804";
		wait for Clk_period;
		Addr <=  "0010011100010";
		Trees_din <= x"ffa414f5";
		wait for Clk_period;
		Addr <=  "0010011100011";
		Trees_din <= x"00a614f5";
		wait for Clk_period;
		Addr <=  "0010011100100";
		Trees_din <= x"3efecf04";
		wait for Clk_period;
		Addr <=  "0010011100101";
		Trees_din <= x"003214f5";
		wait for Clk_period;
		Addr <=  "0010011100110";
		Trees_din <= x"ff6414f5";
		wait for Clk_period;
		Addr <=  "0010011100111";
		Trees_din <= x"81ff3720";
		wait for Clk_period;
		Addr <=  "0010011101000";
		Trees_din <= x"20005e10";
		wait for Clk_period;
		Addr <=  "0010011101001";
		Trees_din <= x"6c003108";
		wait for Clk_period;
		Addr <=  "0010011101010";
		Trees_din <= x"5bfe3a04";
		wait for Clk_period;
		Addr <=  "0010011101011";
		Trees_din <= x"009414f5";
		wait for Clk_period;
		Addr <=  "0010011101100";
		Trees_din <= x"ff8314f5";
		wait for Clk_period;
		Addr <=  "0010011101101";
		Trees_din <= x"2b001d04";
		wait for Clk_period;
		Addr <=  "0010011101110";
		Trees_din <= x"002d14f5";
		wait for Clk_period;
		Addr <=  "0010011101111";
		Trees_din <= x"00d514f5";
		wait for Clk_period;
		Addr <=  "0010011110000";
		Trees_din <= x"5eff9408";
		wait for Clk_period;
		Addr <=  "0010011110001";
		Trees_din <= x"b3fe9604";
		wait for Clk_period;
		Addr <=  "0010011110010";
		Trees_din <= x"ffff14f5";
		wait for Clk_period;
		Addr <=  "0010011110011";
		Trees_din <= x"00c214f5";
		wait for Clk_period;
		Addr <=  "0010011110100";
		Trees_din <= x"0a00d204";
		wait for Clk_period;
		Addr <=  "0010011110101";
		Trees_din <= x"ff7f14f5";
		wait for Clk_period;
		Addr <=  "0010011110110";
		Trees_din <= x"005114f5";
		wait for Clk_period;
		Addr <=  "0010011110111";
		Trees_din <= x"de004310";
		wait for Clk_period;
		Addr <=  "0010011111000";
		Trees_din <= x"efffba08";
		wait for Clk_period;
		Addr <=  "0010011111001";
		Trees_din <= x"edff9904";
		wait for Clk_period;
		Addr <=  "0010011111010";
		Trees_din <= x"fffd14f5";
		wait for Clk_period;
		Addr <=  "0010011111011";
		Trees_din <= x"005114f5";
		wait for Clk_period;
		Addr <=  "0010011111100";
		Trees_din <= x"10002804";
		wait for Clk_period;
		Addr <=  "0010011111101";
		Trees_din <= x"ff9214f5";
		wait for Clk_period;
		Addr <=  "0010011111110";
		Trees_din <= x"001f14f5";
		wait for Clk_period;
		Addr <=  "0010011111111";
		Trees_din <= x"ddfeef08";
		wait for Clk_period;
		Addr <=  "0010100000000";
		Trees_din <= x"a3ffa204";
		wait for Clk_period;
		Addr <=  "0010100000001";
		Trees_din <= x"ffe314f5";
		wait for Clk_period;
		Addr <=  "0010100000010";
		Trees_din <= x"008e14f5";
		wait for Clk_period;
		Addr <=  "0010100000011";
		Trees_din <= x"61002804";
		wait for Clk_period;
		Addr <=  "0010100000100";
		Trees_din <= x"ffa914f5";
		wait for Clk_period;
		Addr <=  "0010100000101";
		Trees_din <= x"005514f5";
		wait for Clk_period;
		Addr <=  "0010100000110";
		Trees_din <= x"c7fe8734";
		wait for Clk_period;
		Addr <=  "0010100000111";
		Trees_din <= x"00ffac20";
		wait for Clk_period;
		Addr <=  "0010100001000";
		Trees_din <= x"2cff2210";
		wait for Clk_period;
		Addr <=  "0010100001001";
		Trees_din <= x"e8ff6d08";
		wait for Clk_period;
		Addr <=  "0010100001010";
		Trees_din <= x"8aff7304";
		wait for Clk_period;
		Addr <=  "0010100001011";
		Trees_din <= x"000414f5";
		wait for Clk_period;
		Addr <=  "0010100001100";
		Trees_din <= x"011414f5";
		wait for Clk_period;
		Addr <=  "0010100001101";
		Trees_din <= x"7a000704";
		wait for Clk_period;
		Addr <=  "0010100001110";
		Trees_din <= x"ff8114f5";
		wait for Clk_period;
		Addr <=  "0010100001111";
		Trees_din <= x"005f14f5";
		wait for Clk_period;
		Addr <=  "0010100010000";
		Trees_din <= x"15000b08";
		wait for Clk_period;
		Addr <=  "0010100010001";
		Trees_din <= x"e8004d04";
		wait for Clk_period;
		Addr <=  "0010100010010";
		Trees_din <= x"ff7314f5";
		wait for Clk_period;
		Addr <=  "0010100010011";
		Trees_din <= x"001714f5";
		wait for Clk_period;
		Addr <=  "0010100010100";
		Trees_din <= x"ceff5a04";
		wait for Clk_period;
		Addr <=  "0010100010101";
		Trees_din <= x"008414f5";
		wait for Clk_period;
		Addr <=  "0010100010110";
		Trees_din <= x"ffcb14f5";
		wait for Clk_period;
		Addr <=  "0010100010111";
		Trees_din <= x"2e000210";
		wait for Clk_period;
		Addr <=  "0010100011000";
		Trees_din <= x"d9ffa508";
		wait for Clk_period;
		Addr <=  "0010100011001";
		Trees_din <= x"95fee804";
		wait for Clk_period;
		Addr <=  "0010100011010";
		Trees_din <= x"ffea14f5";
		wait for Clk_period;
		Addr <=  "0010100011011";
		Trees_din <= x"ff9414f5";
		wait for Clk_period;
		Addr <=  "0010100011100";
		Trees_din <= x"e0ff8204";
		wait for Clk_period;
		Addr <=  "0010100011101";
		Trees_din <= x"009014f5";
		wait for Clk_period;
		Addr <=  "0010100011110";
		Trees_din <= x"ffc414f5";
		wait for Clk_period;
		Addr <=  "0010100011111";
		Trees_din <= x"ff7314f5";
		wait for Clk_period;
		Addr <=  "0010100100000";
		Trees_din <= x"9dffbb20";
		wait for Clk_period;
		Addr <=  "0010100100001";
		Trees_din <= x"7dffe310";
		wait for Clk_period;
		Addr <=  "0010100100010";
		Trees_din <= x"b0ffa208";
		wait for Clk_period;
		Addr <=  "0010100100011";
		Trees_din <= x"e0fea804";
		wait for Clk_period;
		Addr <=  "0010100100100";
		Trees_din <= x"004414f5";
		wait for Clk_period;
		Addr <=  "0010100100101";
		Trees_din <= x"ff7f14f5";
		wait for Clk_period;
		Addr <=  "0010100100110";
		Trees_din <= x"f6feeb04";
		wait for Clk_period;
		Addr <=  "0010100100111";
		Trees_din <= x"ffea14f5";
		wait for Clk_period;
		Addr <=  "0010100101000";
		Trees_din <= x"00cf14f5";
		wait for Clk_period;
		Addr <=  "0010100101001";
		Trees_din <= x"5eff5d08";
		wait for Clk_period;
		Addr <=  "0010100101010";
		Trees_din <= x"77ff3004";
		wait for Clk_period;
		Addr <=  "0010100101011";
		Trees_din <= x"ff7614f5";
		wait for Clk_period;
		Addr <=  "0010100101100";
		Trees_din <= x"fff414f5";
		wait for Clk_period;
		Addr <=  "0010100101101";
		Trees_din <= x"c6ff9204";
		wait for Clk_period;
		Addr <=  "0010100101110";
		Trees_din <= x"006a14f5";
		wait for Clk_period;
		Addr <=  "0010100101111";
		Trees_din <= x"ffc314f5";
		wait for Clk_period;
		Addr <=  "0010100110000";
		Trees_din <= x"50ff040c";
		wait for Clk_period;
		Addr <=  "0010100110001";
		Trees_din <= x"db00d704";
		wait for Clk_period;
		Addr <=  "0010100110010";
		Trees_din <= x"ff6b14f5";
		wait for Clk_period;
		Addr <=  "0010100110011";
		Trees_din <= x"3aff3804";
		wait for Clk_period;
		Addr <=  "0010100110100";
		Trees_din <= x"ffe214f5";
		wait for Clk_period;
		Addr <=  "0010100110101";
		Trees_din <= x"008514f5";
		wait for Clk_period;
		Addr <=  "0010100110110";
		Trees_din <= x"fcfec208";
		wait for Clk_period;
		Addr <=  "0010100110111";
		Trees_din <= x"26008c04";
		wait for Clk_period;
		Addr <=  "0010100111000";
		Trees_din <= x"ff9214f5";
		wait for Clk_period;
		Addr <=  "0010100111001";
		Trees_din <= x"007414f5";
		wait for Clk_period;
		Addr <=  "0010100111010";
		Trees_din <= x"70feef04";
		wait for Clk_period;
		Addr <=  "0010100111011";
		Trees_din <= x"004214f5";
		wait for Clk_period;
		Addr <=  "0010100111100";
		Trees_din <= x"00bb14f5";
		wait for Clk_period;
		Addr <=  "0010100111101";
		Trees_din <= x"eaff4368";
		wait for Clk_period;
		Addr <=  "0010100111110";
		Trees_din <= x"4dfe4d30";
		wait for Clk_period;
		Addr <=  "0010100111111";
		Trees_din <= x"7400171c";
		wait for Clk_period;
		Addr <=  "0010101000000";
		Trees_din <= x"1f00580c";
		wait for Clk_period;
		Addr <=  "0010101000001";
		Trees_din <= x"3effd308";
		wait for Clk_period;
		Addr <=  "0010101000010";
		Trees_din <= x"7ffe6904";
		wait for Clk_period;
		Addr <=  "0010101000011";
		Trees_din <= x"005b1669";
		wait for Clk_period;
		Addr <=  "0010101000100";
		Trees_din <= x"ff671669";
		wait for Clk_period;
		Addr <=  "0010101000101";
		Trees_din <= x"00a31669";
		wait for Clk_period;
		Addr <=  "0010101000110";
		Trees_din <= x"08009e08";
		wait for Clk_period;
		Addr <=  "0010101000111";
		Trees_din <= x"4cfef804";
		wait for Clk_period;
		Addr <=  "0010101001000";
		Trees_din <= x"00dc1669";
		wait for Clk_period;
		Addr <=  "0010101001001";
		Trees_din <= x"00191669";
		wait for Clk_period;
		Addr <=  "0010101001010";
		Trees_din <= x"0a00b204";
		wait for Clk_period;
		Addr <=  "0010101001011";
		Trees_din <= x"ff871669";
		wait for Clk_period;
		Addr <=  "0010101001100";
		Trees_din <= x"003b1669";
		wait for Clk_period;
		Addr <=  "0010101001101";
		Trees_din <= x"36ffac0c";
		wait for Clk_period;
		Addr <=  "0010101001110";
		Trees_din <= x"c9ff7f04";
		wait for Clk_period;
		Addr <=  "0010101001111";
		Trees_din <= x"ffa01669";
		wait for Clk_period;
		Addr <=  "0010101010000";
		Trees_din <= x"c7fe4304";
		wait for Clk_period;
		Addr <=  "0010101010001";
		Trees_din <= x"ffee1669";
		wait for Clk_period;
		Addr <=  "0010101010010";
		Trees_din <= x"00e11669";
		wait for Clk_period;
		Addr <=  "0010101010011";
		Trees_din <= x"a2ff6604";
		wait for Clk_period;
		Addr <=  "0010101010100";
		Trees_din <= x"006d1669";
		wait for Clk_period;
		Addr <=  "0010101010101";
		Trees_din <= x"ff801669";
		wait for Clk_period;
		Addr <=  "0010101010110";
		Trees_din <= x"19fefc1c";
		wait for Clk_period;
		Addr <=  "0010101010111";
		Trees_din <= x"66ffb210";
		wait for Clk_period;
		Addr <=  "0010101011000";
		Trees_din <= x"fcff2308";
		wait for Clk_period;
		Addr <=  "0010101011001";
		Trees_din <= x"e2fea704";
		wait for Clk_period;
		Addr <=  "0010101011010";
		Trees_din <= x"00421669";
		wait for Clk_period;
		Addr <=  "0010101011011";
		Trees_din <= x"01021669";
		wait for Clk_period;
		Addr <=  "0010101011100";
		Trees_din <= x"22011704";
		wait for Clk_period;
		Addr <=  "0010101011101";
		Trees_din <= x"ff981669";
		wait for Clk_period;
		Addr <=  "0010101011110";
		Trees_din <= x"00781669";
		wait for Clk_period;
		Addr <=  "0010101011111";
		Trees_din <= x"1c002608";
		wait for Clk_period;
		Addr <=  "0010101100000";
		Trees_din <= x"21ff6404";
		wait for Clk_period;
		Addr <=  "0010101100001";
		Trees_din <= x"ffee1669";
		wait for Clk_period;
		Addr <=  "0010101100010";
		Trees_din <= x"ff761669";
		wait for Clk_period;
		Addr <=  "0010101100011";
		Trees_din <= x"007c1669";
		wait for Clk_period;
		Addr <=  "0010101100100";
		Trees_din <= x"5100770c";
		wait for Clk_period;
		Addr <=  "0010101100101";
		Trees_din <= x"72ff4004";
		wait for Clk_period;
		Addr <=  "0010101100110";
		Trees_din <= x"008f1669";
		wait for Clk_period;
		Addr <=  "0010101100111";
		Trees_din <= x"00fe7804";
		wait for Clk_period;
		Addr <=  "0010101101000";
		Trees_din <= x"00761669";
		wait for Clk_period;
		Addr <=  "0010101101001";
		Trees_din <= x"ff8e1669";
		wait for Clk_period;
		Addr <=  "0010101101010";
		Trees_din <= x"15ff8408";
		wait for Clk_period;
		Addr <=  "0010101101011";
		Trees_din <= x"ddfed804";
		wait for Clk_period;
		Addr <=  "0010101101100";
		Trees_din <= x"00011669";
		wait for Clk_period;
		Addr <=  "0010101101101";
		Trees_din <= x"ff771669";
		wait for Clk_period;
		Addr <=  "0010101101110";
		Trees_din <= x"c4fea104";
		wait for Clk_period;
		Addr <=  "0010101101111";
		Trees_din <= x"ff8c1669";
		wait for Clk_period;
		Addr <=  "0010101110000";
		Trees_din <= x"00931669";
		wait for Clk_period;
		Addr <=  "0010101110001";
		Trees_din <= x"7eff121c";
		wait for Clk_period;
		Addr <=  "0010101110010";
		Trees_din <= x"d3ffa214";
		wait for Clk_period;
		Addr <=  "0010101110011";
		Trees_din <= x"89fef104";
		wait for Clk_period;
		Addr <=  "0010101110100";
		Trees_din <= x"ff701669";
		wait for Clk_period;
		Addr <=  "0010101110101";
		Trees_din <= x"c7fea708";
		wait for Clk_period;
		Addr <=  "0010101110110";
		Trees_din <= x"3bfef204";
		wait for Clk_period;
		Addr <=  "0010101110111";
		Trees_din <= x"004d1669";
		wait for Clk_period;
		Addr <=  "0010101111000";
		Trees_din <= x"ffde1669";
		wait for Clk_period;
		Addr <=  "0010101111001";
		Trees_din <= x"5a007a04";
		wait for Clk_period;
		Addr <=  "0010101111010";
		Trees_din <= x"00531669";
		wait for Clk_period;
		Addr <=  "0010101111011";
		Trees_din <= x"00111669";
		wait for Clk_period;
		Addr <=  "0010101111100";
		Trees_din <= x"d6ff9b04";
		wait for Clk_period;
		Addr <=  "0010101111101";
		Trees_din <= x"fffe1669";
		wait for Clk_period;
		Addr <=  "0010101111110";
		Trees_din <= x"ff6b1669";
		wait for Clk_period;
		Addr <=  "0010101111111";
		Trees_din <= x"67ffbd1c";
		wait for Clk_period;
		Addr <=  "0010110000000";
		Trees_din <= x"21ff8510";
		wait for Clk_period;
		Addr <=  "0010110000001";
		Trees_din <= x"95ff4608";
		wait for Clk_period;
		Addr <=  "0010110000010";
		Trees_din <= x"1dffa904";
		wait for Clk_period;
		Addr <=  "0010110000011";
		Trees_din <= x"ff6c1669";
		wait for Clk_period;
		Addr <=  "0010110000100";
		Trees_din <= x"00511669";
		wait for Clk_period;
		Addr <=  "0010110000101";
		Trees_din <= x"fcff7104";
		wait for Clk_period;
		Addr <=  "0010110000110";
		Trees_din <= x"009b1669";
		wait for Clk_period;
		Addr <=  "0010110000111";
		Trees_din <= x"ff8a1669";
		wait for Clk_period;
		Addr <=  "0010110001000";
		Trees_din <= x"3700a108";
		wait for Clk_period;
		Addr <=  "0010110001001";
		Trees_din <= x"78003004";
		wait for Clk_period;
		Addr <=  "0010110001010";
		Trees_din <= x"ff801669";
		wait for Clk_period;
		Addr <=  "0010110001011";
		Trees_din <= x"00681669";
		wait for Clk_period;
		Addr <=  "0010110001100";
		Trees_din <= x"00b11669";
		wait for Clk_period;
		Addr <=  "0010110001101";
		Trees_din <= x"1bffc10c";
		wait for Clk_period;
		Addr <=  "0010110001110";
		Trees_din <= x"b9fe9e04";
		wait for Clk_period;
		Addr <=  "0010110001111";
		Trees_din <= x"00a91669";
		wait for Clk_period;
		Addr <=  "0010110010000";
		Trees_din <= x"c7fe5704";
		wait for Clk_period;
		Addr <=  "0010110010001";
		Trees_din <= x"00041669";
		wait for Clk_period;
		Addr <=  "0010110010010";
		Trees_din <= x"ff751669";
		wait for Clk_period;
		Addr <=  "0010110010011";
		Trees_din <= x"b6ff6708";
		wait for Clk_period;
		Addr <=  "0010110010100";
		Trees_din <= x"8dfee804";
		wait for Clk_period;
		Addr <=  "0010110010101";
		Trees_din <= x"013b1669";
		wait for Clk_period;
		Addr <=  "0010110010110";
		Trees_din <= x"00101669";
		wait for Clk_period;
		Addr <=  "0010110010111";
		Trees_din <= x"fdffa004";
		wait for Clk_period;
		Addr <=  "0010110011000";
		Trees_din <= x"ff9c1669";
		wait for Clk_period;
		Addr <=  "0010110011001";
		Trees_din <= x"005f1669";
		wait for Clk_period;
		Addr <=  "0010110011010";
		Trees_din <= x"1aff354c";
		wait for Clk_period;
		Addr <=  "0010110011011";
		Trees_din <= x"bbfff934";
		wait for Clk_period;
		Addr <=  "0010110011100";
		Trees_din <= x"56003620";
		wait for Clk_period;
		Addr <=  "0010110011101";
		Trees_din <= x"6bfe6710";
		wait for Clk_period;
		Addr <=  "0010110011110";
		Trees_din <= x"4dfe3108";
		wait for Clk_period;
		Addr <=  "0010110011111";
		Trees_din <= x"78ff2804";
		wait for Clk_period;
		Addr <=  "0010110100000";
		Trees_din <= x"ffa21765";
		wait for Clk_period;
		Addr <=  "0010110100001";
		Trees_din <= x"006f1765";
		wait for Clk_period;
		Addr <=  "0010110100010";
		Trees_din <= x"56ff0304";
		wait for Clk_period;
		Addr <=  "0010110100011";
		Trees_din <= x"00191765";
		wait for Clk_period;
		Addr <=  "0010110100100";
		Trees_din <= x"ffa01765";
		wait for Clk_period;
		Addr <=  "0010110100101";
		Trees_din <= x"2effee08";
		wait for Clk_period;
		Addr <=  "0010110100110";
		Trees_din <= x"a4ff0d04";
		wait for Clk_period;
		Addr <=  "0010110100111";
		Trees_din <= x"00681765";
		wait for Clk_period;
		Addr <=  "0010110101000";
		Trees_din <= x"000d1765";
		wait for Clk_period;
		Addr <=  "0010110101001";
		Trees_din <= x"52ff3f04";
		wait for Clk_period;
		Addr <=  "0010110101010";
		Trees_din <= x"00201765";
		wait for Clk_period;
		Addr <=  "0010110101011";
		Trees_din <= x"008b1765";
		wait for Clk_period;
		Addr <=  "0010110101100";
		Trees_din <= x"c800890c";
		wait for Clk_period;
		Addr <=  "0010110101101";
		Trees_din <= x"34ffc204";
		wait for Clk_period;
		Addr <=  "0010110101110";
		Trees_din <= x"004a1765";
		wait for Clk_period;
		Addr <=  "0010110101111";
		Trees_din <= x"69fea704";
		wait for Clk_period;
		Addr <=  "0010110110000";
		Trees_din <= x"00441765";
		wait for Clk_period;
		Addr <=  "0010110110001";
		Trees_din <= x"ff691765";
		wait for Clk_period;
		Addr <=  "0010110110010";
		Trees_din <= x"10fef704";
		wait for Clk_period;
		Addr <=  "0010110110011";
		Trees_din <= x"00be1765";
		wait for Clk_period;
		Addr <=  "0010110110100";
		Trees_din <= x"00211765";
		wait for Clk_period;
		Addr <=  "0010110110101";
		Trees_din <= x"a1002614";
		wait for Clk_period;
		Addr <=  "0010110110110";
		Trees_din <= x"3101110c";
		wait for Clk_period;
		Addr <=  "0010110110111";
		Trees_din <= x"eafe8d04";
		wait for Clk_period;
		Addr <=  "0010110111000";
		Trees_din <= x"001f1765";
		wait for Clk_period;
		Addr <=  "0010110111001";
		Trees_din <= x"4dfdbf04";
		wait for Clk_period;
		Addr <=  "0010110111010";
		Trees_din <= x"ffed1765";
		wait for Clk_period;
		Addr <=  "0010110111011";
		Trees_din <= x"ff671765";
		wait for Clk_period;
		Addr <=  "0010110111100";
		Trees_din <= x"94ffa904";
		wait for Clk_period;
		Addr <=  "0010110111101";
		Trees_din <= x"006d1765";
		wait for Clk_period;
		Addr <=  "0010110111110";
		Trees_din <= x"ffcc1765";
		wait for Clk_period;
		Addr <=  "0010110111111";
		Trees_din <= x"007c1765";
		wait for Clk_period;
		Addr <=  "0010111000000";
		Trees_din <= x"1bff790c";
		wait for Clk_period;
		Addr <=  "0010111000001";
		Trees_din <= x"8800ae08";
		wait for Clk_period;
		Addr <=  "0010111000010";
		Trees_din <= x"f0fe3604";
		wait for Clk_period;
		Addr <=  "0010111000011";
		Trees_din <= x"00261765";
		wait for Clk_period;
		Addr <=  "0010111000100";
		Trees_din <= x"ff661765";
		wait for Clk_period;
		Addr <=  "0010111000101";
		Trees_din <= x"00571765";
		wait for Clk_period;
		Addr <=  "0010111000110";
		Trees_din <= x"18003d1c";
		wait for Clk_period;
		Addr <=  "0010111000111";
		Trees_din <= x"da008810";
		wait for Clk_period;
		Addr <=  "0010111001000";
		Trees_din <= x"17002b08";
		wait for Clk_period;
		Addr <=  "0010111001001";
		Trees_din <= x"b8ff4804";
		wait for Clk_period;
		Addr <=  "0010111001010";
		Trees_din <= x"003f1765";
		wait for Clk_period;
		Addr <=  "0010111001011";
		Trees_din <= x"ff9d1765";
		wait for Clk_period;
		Addr <=  "0010111001100";
		Trees_din <= x"a7ff7d04";
		wait for Clk_period;
		Addr <=  "0010111001101";
		Trees_din <= x"ffb41765";
		wait for Clk_period;
		Addr <=  "0010111001110";
		Trees_din <= x"00a21765";
		wait for Clk_period;
		Addr <=  "0010111001111";
		Trees_din <= x"4cff6108";
		wait for Clk_period;
		Addr <=  "0010111010000";
		Trees_din <= x"e4ff0704";
		wait for Clk_period;
		Addr <=  "0010111010001";
		Trees_din <= x"00f31765";
		wait for Clk_period;
		Addr <=  "0010111010010";
		Trees_din <= x"00171765";
		wait for Clk_period;
		Addr <=  "0010111010011";
		Trees_din <= x"ffe01765";
		wait for Clk_period;
		Addr <=  "0010111010100";
		Trees_din <= x"44ff6e04";
		wait for Clk_period;
		Addr <=  "0010111010101";
		Trees_din <= x"008c1765";
		wait for Clk_period;
		Addr <=  "0010111010110";
		Trees_din <= x"4efff404";
		wait for Clk_period;
		Addr <=  "0010111010111";
		Trees_din <= x"ff691765";
		wait for Clk_period;
		Addr <=  "0010111011000";
		Trees_din <= x"00191765";
		wait for Clk_period;
		Addr <=  "0010111011001";
		Trees_din <= x"19ffa044";
		wait for Clk_period;
		Addr <=  "0010111011010";
		Trees_din <= x"6f003e34";
		wait for Clk_period;
		Addr <=  "0010111011011";
		Trees_din <= x"81fef514";
		wait for Clk_period;
		Addr <=  "0010111011100";
		Trees_din <= x"8affe704";
		wait for Clk_period;
		Addr <=  "0010111011101";
		Trees_din <= x"ff681869";
		wait for Clk_period;
		Addr <=  "0010111011110";
		Trees_din <= x"2effab08";
		wait for Clk_period;
		Addr <=  "0010111011111";
		Trees_din <= x"2dff9304";
		wait for Clk_period;
		Addr <=  "0010111100000";
		Trees_din <= x"00981869";
		wait for Clk_period;
		Addr <=  "0010111100001";
		Trees_din <= x"ffa71869";
		wait for Clk_period;
		Addr <=  "0010111100010";
		Trees_din <= x"f7ff8704";
		wait for Clk_period;
		Addr <=  "0010111100011";
		Trees_din <= x"ff831869";
		wait for Clk_period;
		Addr <=  "0010111100100";
		Trees_din <= x"ffe41869";
		wait for Clk_period;
		Addr <=  "0010111100101";
		Trees_din <= x"90ff5110";
		wait for Clk_period;
		Addr <=  "0010111100110";
		Trees_din <= x"dcffb708";
		wait for Clk_period;
		Addr <=  "0010111100111";
		Trees_din <= x"70ff2904";
		wait for Clk_period;
		Addr <=  "0010111101000";
		Trees_din <= x"00011869";
		wait for Clk_period;
		Addr <=  "0010111101001";
		Trees_din <= x"00761869";
		wait for Clk_period;
		Addr <=  "0010111101010";
		Trees_din <= x"82ffaa04";
		wait for Clk_period;
		Addr <=  "0010111101011";
		Trees_din <= x"ffb61869";
		wait for Clk_period;
		Addr <=  "0010111101100";
		Trees_din <= x"00201869";
		wait for Clk_period;
		Addr <=  "0010111101101";
		Trees_din <= x"8ffe5708";
		wait for Clk_period;
		Addr <=  "0010111101110";
		Trees_din <= x"eeffe704";
		wait for Clk_period;
		Addr <=  "0010111101111";
		Trees_din <= x"00041869";
		wait for Clk_period;
		Addr <=  "0010111110000";
		Trees_din <= x"00c41869";
		wait for Clk_period;
		Addr <=  "0010111110001";
		Trees_din <= x"a2ffd204";
		wait for Clk_period;
		Addr <=  "0010111110010";
		Trees_din <= x"00331869";
		wait for Clk_period;
		Addr <=  "0010111110011";
		Trees_din <= x"fffc1869";
		wait for Clk_period;
		Addr <=  "0010111110100";
		Trees_din <= x"3eff1a08";
		wait for Clk_period;
		Addr <=  "0010111110101";
		Trees_din <= x"d600eb04";
		wait for Clk_period;
		Addr <=  "0010111110110";
		Trees_din <= x"ffeb1869";
		wait for Clk_period;
		Addr <=  "0010111110111";
		Trees_din <= x"009b1869";
		wait for Clk_period;
		Addr <=  "0010111111000";
		Trees_din <= x"c1ffb104";
		wait for Clk_period;
		Addr <=  "0010111111001";
		Trees_din <= x"ff681869";
		wait for Clk_period;
		Addr <=  "0010111111010";
		Trees_din <= x"00051869";
		wait for Clk_period;
		Addr <=  "0010111111011";
		Trees_din <= x"db00ac20";
		wait for Clk_period;
		Addr <=  "0010111111100";
		Trees_din <= x"dc007a10";
		wait for Clk_period;
		Addr <=  "0010111111101";
		Trees_din <= x"4400b408";
		wait for Clk_period;
		Addr <=  "0010111111110";
		Trees_din <= x"dffe8104";
		wait for Clk_period;
		Addr <=  "0010111111111";
		Trees_din <= x"00381869";
		wait for Clk_period;
		Addr <=  "0011000000000";
		Trees_din <= x"ff651869";
		wait for Clk_period;
		Addr <=  "0011000000001";
		Trees_din <= x"1fffe004";
		wait for Clk_period;
		Addr <=  "0011000000010";
		Trees_din <= x"ffe61869";
		wait for Clk_period;
		Addr <=  "0011000000011";
		Trees_din <= x"005c1869";
		wait for Clk_period;
		Addr <=  "0011000000100";
		Trees_din <= x"67ff5604";
		wait for Clk_period;
		Addr <=  "0011000000101";
		Trees_din <= x"ff981869";
		wait for Clk_period;
		Addr <=  "0011000000110";
		Trees_din <= x"d7009608";
		wait for Clk_period;
		Addr <=  "0011000000111";
		Trees_din <= x"d0006404";
		wait for Clk_period;
		Addr <=  "0011000001000";
		Trees_din <= x"00b51869";
		wait for Clk_period;
		Addr <=  "0011000001001";
		Trees_din <= x"00321869";
		wait for Clk_period;
		Addr <=  "0011000001010";
		Trees_din <= x"ffd71869";
		wait for Clk_period;
		Addr <=  "0011000001011";
		Trees_din <= x"e0fef308";
		wait for Clk_period;
		Addr <=  "0011000001100";
		Trees_din <= x"4dfebb04";
		wait for Clk_period;
		Addr <=  "0011000001101";
		Trees_din <= x"ff8b1869";
		wait for Clk_period;
		Addr <=  "0011000001110";
		Trees_din <= x"ffe11869";
		wait for Clk_period;
		Addr <=  "0011000001111";
		Trees_din <= x"b1fecc08";
		wait for Clk_period;
		Addr <=  "0011000010000";
		Trees_din <= x"aaff3804";
		wait for Clk_period;
		Addr <=  "0011000010001";
		Trees_din <= x"00d31869";
		wait for Clk_period;
		Addr <=  "0011000010010";
		Trees_din <= x"002d1869";
		wait for Clk_period;
		Addr <=  "0011000010011";
		Trees_din <= x"99ff3908";
		wait for Clk_period;
		Addr <=  "0011000010100";
		Trees_din <= x"acffe504";
		wait for Clk_period;
		Addr <=  "0011000010101";
		Trees_din <= x"fffe1869";
		wait for Clk_period;
		Addr <=  "0011000010110";
		Trees_din <= x"ff8a1869";
		wait for Clk_period;
		Addr <=  "0011000010111";
		Trees_din <= x"d2fec404";
		wait for Clk_period;
		Addr <=  "0011000011000";
		Trees_din <= x"00a71869";
		wait for Clk_period;
		Addr <=  "0011000011001";
		Trees_din <= x"fff01869";
		wait for Clk_period;
		Addr <=  "0011000011010";
		Trees_din <= x"89008268";
		wait for Clk_period;
		Addr <=  "0011000011011";
		Trees_din <= x"9dff4e28";
		wait for Clk_period;
		Addr <=  "0011000011100";
		Trees_din <= x"f0003620";
		wait for Clk_period;
		Addr <=  "0011000011101";
		Trees_din <= x"8aff5010";
		wait for Clk_period;
		Addr <=  "0011000011110";
		Trees_din <= x"94ff9f08";
		wait for Clk_period;
		Addr <=  "0011000011111";
		Trees_din <= x"34004104";
		wait for Clk_period;
		Addr <=  "0011000100000";
		Trees_din <= x"ff7919a5";
		wait for Clk_period;
		Addr <=  "0011000100001";
		Trees_din <= x"001119a5";
		wait for Clk_period;
		Addr <=  "0011000100010";
		Trees_din <= x"53ff2104";
		wait for Clk_period;
		Addr <=  "0011000100011";
		Trees_din <= x"ff8519a5";
		wait for Clk_period;
		Addr <=  "0011000100100";
		Trees_din <= x"007419a5";
		wait for Clk_period;
		Addr <=  "0011000100101";
		Trees_din <= x"b9fe4008";
		wait for Clk_period;
		Addr <=  "0011000100110";
		Trees_din <= x"6cffe904";
		wait for Clk_period;
		Addr <=  "0011000100111";
		Trees_din <= x"ffd219a5";
		wait for Clk_period;
		Addr <=  "0011000101000";
		Trees_din <= x"00b119a5";
		wait for Clk_period;
		Addr <=  "0011000101001";
		Trees_din <= x"b3ffbd04";
		wait for Clk_period;
		Addr <=  "0011000101010";
		Trees_din <= x"ff8f19a5";
		wait for Clk_period;
		Addr <=  "0011000101011";
		Trees_din <= x"003b19a5";
		wait for Clk_period;
		Addr <=  "0011000101100";
		Trees_din <= x"57ff0f04";
		wait for Clk_period;
		Addr <=  "0011000101101";
		Trees_din <= x"00d419a5";
		wait for Clk_period;
		Addr <=  "0011000101110";
		Trees_din <= x"ffe419a5";
		wait for Clk_period;
		Addr <=  "0011000101111";
		Trees_din <= x"ab007120";
		wait for Clk_period;
		Addr <=  "0011000110000";
		Trees_din <= x"24ffdc10";
		wait for Clk_period;
		Addr <=  "0011000110001";
		Trees_din <= x"2b004208";
		wait for Clk_period;
		Addr <=  "0011000110010";
		Trees_din <= x"0bffa504";
		wait for Clk_period;
		Addr <=  "0011000110011";
		Trees_din <= x"ff7719a5";
		wait for Clk_period;
		Addr <=  "0011000110100";
		Trees_din <= x"ffdc19a5";
		wait for Clk_period;
		Addr <=  "0011000110101";
		Trees_din <= x"b3ff3504";
		wait for Clk_period;
		Addr <=  "0011000110110";
		Trees_din <= x"ffbd19a5";
		wait for Clk_period;
		Addr <=  "0011000110111";
		Trees_din <= x"009719a5";
		wait for Clk_period;
		Addr <=  "0011000111000";
		Trees_din <= x"2dfeba08";
		wait for Clk_period;
		Addr <=  "0011000111001";
		Trees_din <= x"b2ffe704";
		wait for Clk_period;
		Addr <=  "0011000111010";
		Trees_din <= x"00af19a5";
		wait for Clk_period;
		Addr <=  "0011000111011";
		Trees_din <= x"ffe819a5";
		wait for Clk_period;
		Addr <=  "0011000111100";
		Trees_din <= x"a2ffdd04";
		wait for Clk_period;
		Addr <=  "0011000111101";
		Trees_din <= x"002919a5";
		wait for Clk_period;
		Addr <=  "0011000111110";
		Trees_din <= x"ff9e19a5";
		wait for Clk_period;
		Addr <=  "0011000111111";
		Trees_din <= x"c7fe7910";
		wait for Clk_period;
		Addr <=  "0011001000000";
		Trees_din <= x"ebff3508";
		wait for Clk_period;
		Addr <=  "0011001000001";
		Trees_din <= x"4bff4704";
		wait for Clk_period;
		Addr <=  "0011001000010";
		Trees_din <= x"ff9819a5";
		wait for Clk_period;
		Addr <=  "0011001000011";
		Trees_din <= x"003619a5";
		wait for Clk_period;
		Addr <=  "0011001000100";
		Trees_din <= x"41ff3f04";
		wait for Clk_period;
		Addr <=  "0011001000101";
		Trees_din <= x"fffa19a5";
		wait for Clk_period;
		Addr <=  "0011001000110";
		Trees_din <= x"00a919a5";
		wait for Clk_period;
		Addr <=  "0011001000111";
		Trees_din <= x"1dfe9f08";
		wait for Clk_period;
		Addr <=  "0011001001000";
		Trees_din <= x"4eff9f04";
		wait for Clk_period;
		Addr <=  "0011001001001";
		Trees_din <= x"ff7b19a5";
		wait for Clk_period;
		Addr <=  "0011001001010";
		Trees_din <= x"003719a5";
		wait for Clk_period;
		Addr <=  "0011001001011";
		Trees_din <= x"b8ffa604";
		wait for Clk_period;
		Addr <=  "0011001001100";
		Trees_din <= x"005d19a5";
		wait for Clk_period;
		Addr <=  "0011001001101";
		Trees_din <= x"000e19a5";
		wait for Clk_period;
		Addr <=  "0011001001110";
		Trees_din <= x"a4ffdb28";
		wait for Clk_period;
		Addr <=  "0011001001111";
		Trees_din <= x"19ff821c";
		wait for Clk_period;
		Addr <=  "0011001010000";
		Trees_din <= x"84ff520c";
		wait for Clk_period;
		Addr <=  "0011001010001";
		Trees_din <= x"4dfebe04";
		wait for Clk_period;
		Addr <=  "0011001010010";
		Trees_din <= x"ff7619a5";
		wait for Clk_period;
		Addr <=  "0011001010011";
		Trees_din <= x"87ff8604";
		wait for Clk_period;
		Addr <=  "0011001010100";
		Trees_din <= x"ffae19a5";
		wait for Clk_period;
		Addr <=  "0011001010101";
		Trees_din <= x"00bf19a5";
		wait for Clk_period;
		Addr <=  "0011001010110";
		Trees_din <= x"61ffac08";
		wait for Clk_period;
		Addr <=  "0011001010111";
		Trees_din <= x"4dfeb904";
		wait for Clk_period;
		Addr <=  "0011001011000";
		Trees_din <= x"009519a5";
		wait for Clk_period;
		Addr <=  "0011001011001";
		Trees_din <= x"000719a5";
		wait for Clk_period;
		Addr <=  "0011001011010";
		Trees_din <= x"cdffec04";
		wait for Clk_period;
		Addr <=  "0011001011011";
		Trees_din <= x"ff7719a5";
		wait for Clk_period;
		Addr <=  "0011001011100";
		Trees_din <= x"005519a5";
		wait for Clk_period;
		Addr <=  "0011001011101";
		Trees_din <= x"15006308";
		wait for Clk_period;
		Addr <=  "0011001011110";
		Trees_din <= x"a5ff7204";
		wait for Clk_period;
		Addr <=  "0011001011111";
		Trees_din <= x"ff7219a5";
		wait for Clk_period;
		Addr <=  "0011001100000";
		Trees_din <= x"000b19a5";
		wait for Clk_period;
		Addr <=  "0011001100001";
		Trees_din <= x"006319a5";
		wait for Clk_period;
		Addr <=  "0011001100010";
		Trees_din <= x"20007c08";
		wait for Clk_period;
		Addr <=  "0011001100011";
		Trees_din <= x"5eff8804";
		wait for Clk_period;
		Addr <=  "0011001100100";
		Trees_din <= x"ffef19a5";
		wait for Clk_period;
		Addr <=  "0011001100101";
		Trees_din <= x"ff7019a5";
		wait for Clk_period;
		Addr <=  "0011001100110";
		Trees_din <= x"4dfde104";
		wait for Clk_period;
		Addr <=  "0011001100111";
		Trees_din <= x"007519a5";
		wait for Clk_period;
		Addr <=  "0011001101000";
		Trees_din <= x"ffda19a5";
		wait for Clk_period;
		Addr <=  "0011001101001";
		Trees_din <= x"fcfebc38";
		wait for Clk_period;
		Addr <=  "0011001101010";
		Trees_din <= x"1fffba0c";
		wait for Clk_period;
		Addr <=  "0011001101011";
		Trees_din <= x"0b006304";
		wait for Clk_period;
		Addr <=  "0011001101100";
		Trees_din <= x"ff6a1b09";
		wait for Clk_period;
		Addr <=  "0011001101101";
		Trees_din <= x"f0ff6804";
		wait for Clk_period;
		Addr <=  "0011001101110";
		Trees_din <= x"ffa21b09";
		wait for Clk_period;
		Addr <=  "0011001101111";
		Trees_din <= x"006a1b09";
		wait for Clk_period;
		Addr <=  "0011001110000";
		Trees_din <= x"fbff8814";
		wait for Clk_period;
		Addr <=  "0011001110001";
		Trees_din <= x"f202a008";
		wait for Clk_period;
		Addr <=  "0011001110010";
		Trees_din <= x"2cff5304";
		wait for Clk_period;
		Addr <=  "0011001110011";
		Trees_din <= x"005c1b09";
		wait for Clk_period;
		Addr <=  "0011001110100";
		Trees_din <= x"ff8e1b09";
		wait for Clk_period;
		Addr <=  "0011001110101";
		Trees_din <= x"d2fe9e08";
		wait for Clk_period;
		Addr <=  "0011001110110";
		Trees_din <= x"bfffaa04";
		wait for Clk_period;
		Addr <=  "0011001110111";
		Trees_din <= x"00bc1b09";
		wait for Clk_period;
		Addr <=  "0011001111000";
		Trees_din <= x"00271b09";
		wait for Clk_period;
		Addr <=  "0011001111001";
		Trees_din <= x"ffd51b09";
		wait for Clk_period;
		Addr <=  "0011001111010";
		Trees_din <= x"74ffc50c";
		wait for Clk_period;
		Addr <=  "0011001111011";
		Trees_din <= x"e2ff4204";
		wait for Clk_period;
		Addr <=  "0011001111100";
		Trees_din <= x"ffae1b09";
		wait for Clk_period;
		Addr <=  "0011001111101";
		Trees_din <= x"36ffaa04";
		wait for Clk_period;
		Addr <=  "0011001111110";
		Trees_din <= x"00351b09";
		wait for Clk_period;
		Addr <=  "0011001111111";
		Trees_din <= x"00b21b09";
		wait for Clk_period;
		Addr <=  "0011010000000";
		Trees_din <= x"69fee808";
		wait for Clk_period;
		Addr <=  "0011010000001";
		Trees_din <= x"7d000104";
		wait for Clk_period;
		Addr <=  "0011010000010";
		Trees_din <= x"ffb01b09";
		wait for Clk_period;
		Addr <=  "0011010000011";
		Trees_din <= x"005a1b09";
		wait for Clk_period;
		Addr <=  "0011010000100";
		Trees_din <= x"ff6b1b09";
		wait for Clk_period;
		Addr <=  "0011010000101";
		Trees_din <= x"b4ff3b40";
		wait for Clk_period;
		Addr <=  "0011010000110";
		Trees_din <= x"a3ff3020";
		wait for Clk_period;
		Addr <=  "0011010000111";
		Trees_din <= x"49ff8f10";
		wait for Clk_period;
		Addr <=  "0011010001000";
		Trees_din <= x"d6006b08";
		wait for Clk_period;
		Addr <=  "0011010001001";
		Trees_din <= x"2c001104";
		wait for Clk_period;
		Addr <=  "0011010001010";
		Trees_din <= x"ff851b09";
		wait for Clk_period;
		Addr <=  "0011010001011";
		Trees_din <= x"00391b09";
		wait for Clk_period;
		Addr <=  "0011010001100";
		Trees_din <= x"b0ff1204";
		wait for Clk_period;
		Addr <=  "0011010001101";
		Trees_din <= x"ffa81b09";
		wait for Clk_period;
		Addr <=  "0011010001110";
		Trees_din <= x"00be1b09";
		wait for Clk_period;
		Addr <=  "0011010001111";
		Trees_din <= x"1b00a208";
		wait for Clk_period;
		Addr <=  "0011010010000";
		Trees_din <= x"53ff9504";
		wait for Clk_period;
		Addr <=  "0011010010001";
		Trees_din <= x"ffee1b09";
		wait for Clk_period;
		Addr <=  "0011010010010";
		Trees_din <= x"ff811b09";
		wait for Clk_period;
		Addr <=  "0011010010011";
		Trees_din <= x"8efffb04";
		wait for Clk_period;
		Addr <=  "0011010010100";
		Trees_din <= x"008a1b09";
		wait for Clk_period;
		Addr <=  "0011010010101";
		Trees_din <= x"ffad1b09";
		wait for Clk_period;
		Addr <=  "0011010010110";
		Trees_din <= x"beffbb10";
		wait for Clk_period;
		Addr <=  "0011010010111";
		Trees_din <= x"9dffc108";
		wait for Clk_period;
		Addr <=  "0011010011000";
		Trees_din <= x"acfffa04";
		wait for Clk_period;
		Addr <=  "0011010011001";
		Trees_din <= x"001b1b09";
		wait for Clk_period;
		Addr <=  "0011010011010";
		Trees_din <= x"ff9a1b09";
		wait for Clk_period;
		Addr <=  "0011010011011";
		Trees_din <= x"9cff9a04";
		wait for Clk_period;
		Addr <=  "0011010011100";
		Trees_din <= x"005e1b09";
		wait for Clk_period;
		Addr <=  "0011010011101";
		Trees_din <= x"ffcb1b09";
		wait for Clk_period;
		Addr <=  "0011010011110";
		Trees_din <= x"80ff5808";
		wait for Clk_period;
		Addr <=  "0011010011111";
		Trees_din <= x"1cff4904";
		wait for Clk_period;
		Addr <=  "0011010100000";
		Trees_din <= x"ffb51b09";
		wait for Clk_period;
		Addr <=  "0011010100001";
		Trees_din <= x"00311b09";
		wait for Clk_period;
		Addr <=  "0011010100010";
		Trees_din <= x"45feec04";
		wait for Clk_period;
		Addr <=  "0011010100011";
		Trees_din <= x"002c1b09";
		wait for Clk_period;
		Addr <=  "0011010100100";
		Trees_din <= x"00781b09";
		wait for Clk_period;
		Addr <=  "0011010100101";
		Trees_din <= x"70ff2720";
		wait for Clk_period;
		Addr <=  "0011010100110";
		Trees_din <= x"9bff1110";
		wait for Clk_period;
		Addr <=  "0011010100111";
		Trees_din <= x"b7ff4a08";
		wait for Clk_period;
		Addr <=  "0011010101000";
		Trees_din <= x"2200bf04";
		wait for Clk_period;
		Addr <=  "0011010101001";
		Trees_din <= x"ff9c1b09";
		wait for Clk_period;
		Addr <=  "0011010101010";
		Trees_din <= x"005d1b09";
		wait for Clk_period;
		Addr <=  "0011010101011";
		Trees_din <= x"2bfee304";
		wait for Clk_period;
		Addr <=  "0011010101100";
		Trees_din <= x"00341b09";
		wait for Clk_period;
		Addr <=  "0011010101101";
		Trees_din <= x"ff621b09";
		wait for Clk_period;
		Addr <=  "0011010101110";
		Trees_din <= x"86ff7608";
		wait for Clk_period;
		Addr <=  "0011010101111";
		Trees_din <= x"2effa904";
		wait for Clk_period;
		Addr <=  "0011010110000";
		Trees_din <= x"ff931b09";
		wait for Clk_period;
		Addr <=  "0011010110001";
		Trees_din <= x"000f1b09";
		wait for Clk_period;
		Addr <=  "0011010110010";
		Trees_din <= x"36fef704";
		wait for Clk_period;
		Addr <=  "0011010110011";
		Trees_din <= x"ff801b09";
		wait for Clk_period;
		Addr <=  "0011010110100";
		Trees_din <= x"00681b09";
		wait for Clk_period;
		Addr <=  "0011010110101";
		Trees_din <= x"28fee60c";
		wait for Clk_period;
		Addr <=  "0011010110110";
		Trees_din <= x"38ff2404";
		wait for Clk_period;
		Addr <=  "0011010110111";
		Trees_din <= x"ff961b09";
		wait for Clk_period;
		Addr <=  "0011010111000";
		Trees_din <= x"4aff5c04";
		wait for Clk_period;
		Addr <=  "0011010111001";
		Trees_din <= x"00cf1b09";
		wait for Clk_period;
		Addr <=  "0011010111010";
		Trees_din <= x"ffcf1b09";
		wait for Clk_period;
		Addr <=  "0011010111011";
		Trees_din <= x"d000bb08";
		wait for Clk_period;
		Addr <=  "0011010111100";
		Trees_din <= x"d4fefd04";
		wait for Clk_period;
		Addr <=  "0011010111101";
		Trees_din <= x"00681b09";
		wait for Clk_period;
		Addr <=  "0011010111110";
		Trees_din <= x"ffbb1b09";
		wait for Clk_period;
		Addr <=  "0011010111111";
		Trees_din <= x"d5ffe604";
		wait for Clk_period;
		Addr <=  "0011011000000";
		Trees_din <= x"ffbd1b09";
		wait for Clk_period;
		Addr <=  "0011011000001";
		Trees_din <= x"00b61b09";
		wait for Clk_period;
		Addr <=  "0011011000010";
		Trees_din <= x"1aff3554";
		wait for Clk_period;
		Addr <=  "0011011000011";
		Trees_din <= x"bbfff940";
		wait for Clk_period;
		Addr <=  "0011011000100";
		Trees_din <= x"61fece20";
		wait for Clk_period;
		Addr <=  "0011011000101";
		Trees_din <= x"31000210";
		wait for Clk_period;
		Addr <=  "0011011000110";
		Trees_din <= x"09006408";
		wait for Clk_period;
		Addr <=  "0011011000111";
		Trees_din <= x"a6001304";
		wait for Clk_period;
		Addr <=  "0011011001000";
		Trees_din <= x"ff761c1d";
		wait for Clk_period;
		Addr <=  "0011011001001";
		Trees_din <= x"00291c1d";
		wait for Clk_period;
		Addr <=  "0011011001010";
		Trees_din <= x"72004304";
		wait for Clk_period;
		Addr <=  "0011011001011";
		Trees_din <= x"000b1c1d";
		wait for Clk_period;
		Addr <=  "0011011001100";
		Trees_din <= x"00701c1d";
		wait for Clk_period;
		Addr <=  "0011011001101";
		Trees_din <= x"4dfe5008";
		wait for Clk_period;
		Addr <=  "0011011001110";
		Trees_din <= x"0cfebf04";
		wait for Clk_period;
		Addr <=  "0011011001111";
		Trees_din <= x"ffe21c1d";
		wait for Clk_period;
		Addr <=  "0011011010000";
		Trees_din <= x"009b1c1d";
		wait for Clk_period;
		Addr <=  "0011011010001";
		Trees_din <= x"8eff9d04";
		wait for Clk_period;
		Addr <=  "0011011010010";
		Trees_din <= x"00571c1d";
		wait for Clk_period;
		Addr <=  "0011011010011";
		Trees_din <= x"ffb11c1d";
		wait for Clk_period;
		Addr <=  "0011011010100";
		Trees_din <= x"91002710";
		wait for Clk_period;
		Addr <=  "0011011010101";
		Trees_din <= x"faff7808";
		wait for Clk_period;
		Addr <=  "0011011010110";
		Trees_din <= x"2bffdf04";
		wait for Clk_period;
		Addr <=  "0011011010111";
		Trees_din <= x"00141c1d";
		wait for Clk_period;
		Addr <=  "0011011011000";
		Trees_din <= x"00581c1d";
		wait for Clk_period;
		Addr <=  "0011011011001";
		Trees_din <= x"db00c404";
		wait for Clk_period;
		Addr <=  "0011011011010";
		Trees_din <= x"fff31c1d";
		wait for Clk_period;
		Addr <=  "0011011011011";
		Trees_din <= x"00491c1d";
		wait for Clk_period;
		Addr <=  "0011011011100";
		Trees_din <= x"0fff1808";
		wait for Clk_period;
		Addr <=  "0011011011101";
		Trees_din <= x"b4febc04";
		wait for Clk_period;
		Addr <=  "0011011011110";
		Trees_din <= x"00721c1d";
		wait for Clk_period;
		Addr <=  "0011011011111";
		Trees_din <= x"ffc81c1d";
		wait for Clk_period;
		Addr <=  "0011011100000";
		Trees_din <= x"58fe6904";
		wait for Clk_period;
		Addr <=  "0011011100001";
		Trees_din <= x"fff01c1d";
		wait for Clk_period;
		Addr <=  "0011011100010";
		Trees_din <= x"ff701c1d";
		wait for Clk_period;
		Addr <=  "0011011100011";
		Trees_din <= x"a1002610";
		wait for Clk_period;
		Addr <=  "0011011100100";
		Trees_din <= x"3101110c";
		wait for Clk_period;
		Addr <=  "0011011100101";
		Trees_din <= x"eafe8d04";
		wait for Clk_period;
		Addr <=  "0011011100110";
		Trees_din <= x"001f1c1d";
		wait for Clk_period;
		Addr <=  "0011011100111";
		Trees_din <= x"4dfdbf04";
		wait for Clk_period;
		Addr <=  "0011011101000";
		Trees_din <= x"ffed1c1d";
		wait for Clk_period;
		Addr <=  "0011011101001";
		Trees_din <= x"ff6c1c1d";
		wait for Clk_period;
		Addr <=  "0011011101010";
		Trees_din <= x"002e1c1d";
		wait for Clk_period;
		Addr <=  "0011011101011";
		Trees_din <= x"00661c1d";
		wait for Clk_period;
		Addr <=  "0011011101100";
		Trees_din <= x"1bff790c";
		wait for Clk_period;
		Addr <=  "0011011101101";
		Trees_din <= x"8800ae08";
		wait for Clk_period;
		Addr <=  "0011011101110";
		Trees_din <= x"b9fe6f04";
		wait for Clk_period;
		Addr <=  "0011011101111";
		Trees_din <= x"00131c1d";
		wait for Clk_period;
		Addr <=  "0011011110000";
		Trees_din <= x"ff6a1c1d";
		wait for Clk_period;
		Addr <=  "0011011110001";
		Trees_din <= x"00491c1d";
		wait for Clk_period;
		Addr <=  "0011011110010";
		Trees_din <= x"cfff8e10";
		wait for Clk_period;
		Addr <=  "0011011110011";
		Trees_din <= x"92ff0d04";
		wait for Clk_period;
		Addr <=  "0011011110100";
		Trees_din <= x"ff9d1c1d";
		wait for Clk_period;
		Addr <=  "0011011110101";
		Trees_din <= x"fcff0404";
		wait for Clk_period;
		Addr <=  "0011011110110";
		Trees_din <= x"00041c1d";
		wait for Clk_period;
		Addr <=  "0011011110111";
		Trees_din <= x"9cff7804";
		wait for Clk_period;
		Addr <=  "0011011111000";
		Trees_din <= x"010d1c1d";
		wait for Clk_period;
		Addr <=  "0011011111001";
		Trees_din <= x"003f1c1d";
		wait for Clk_period;
		Addr <=  "0011011111010";
		Trees_din <= x"39ffa110";
		wait for Clk_period;
		Addr <=  "0011011111011";
		Trees_din <= x"feff8108";
		wait for Clk_period;
		Addr <=  "0011011111100";
		Trees_din <= x"70ff0e04";
		wait for Clk_period;
		Addr <=  "0011011111101";
		Trees_din <= x"fff01c1d";
		wait for Clk_period;
		Addr <=  "0011011111110";
		Trees_din <= x"00ae1c1d";
		wait for Clk_period;
		Addr <=  "0011011111111";
		Trees_din <= x"1cffab04";
		wait for Clk_period;
		Addr <=  "0011100000000";
		Trees_din <= x"ff961c1d";
		wait for Clk_period;
		Addr <=  "0011100000001";
		Trees_din <= x"00561c1d";
		wait for Clk_period;
		Addr <=  "0011100000010";
		Trees_din <= x"a5fe8e04";
		wait for Clk_period;
		Addr <=  "0011100000011";
		Trees_din <= x"00831c1d";
		wait for Clk_period;
		Addr <=  "0011100000100";
		Trees_din <= x"88009504";
		wait for Clk_period;
		Addr <=  "0011100000101";
		Trees_din <= x"ff741c1d";
		wait for Clk_period;
		Addr <=  "0011100000110";
		Trees_din <= x"002d1c1d";
		wait for Clk_period;
		Addr <=  "0011100000111";
		Trees_din <= x"19ffa05c";
		wait for Clk_period;
		Addr <=  "0011100001000";
		Trees_din <= x"20feec1c";
		wait for Clk_period;
		Addr <=  "0011100001001";
		Trees_din <= x"35fe8d10";
		wait for Clk_period;
		Addr <=  "0011100001010";
		Trees_din <= x"e4fe9304";
		wait for Clk_period;
		Addr <=  "0011100001011";
		Trees_din <= x"ff8d1d39";
		wait for Clk_period;
		Addr <=  "0011100001100";
		Trees_din <= x"35fe5e04";
		wait for Clk_period;
		Addr <=  "0011100001101";
		Trees_din <= x"ffde1d39";
		wait for Clk_period;
		Addr <=  "0011100001110";
		Trees_din <= x"1afed304";
		wait for Clk_period;
		Addr <=  "0011100001111";
		Trees_din <= x"00bf1d39";
		wait for Clk_period;
		Addr <=  "0011100010000";
		Trees_din <= x"00241d39";
		wait for Clk_period;
		Addr <=  "0011100010001";
		Trees_din <= x"a5fe8004";
		wait for Clk_period;
		Addr <=  "0011100010010";
		Trees_din <= x"004e1d39";
		wait for Clk_period;
		Addr <=  "0011100010011";
		Trees_din <= x"2dffb704";
		wait for Clk_period;
		Addr <=  "0011100010100";
		Trees_din <= x"ff6a1d39";
		wait for Clk_period;
		Addr <=  "0011100010101";
		Trees_din <= x"00291d39";
		wait for Clk_period;
		Addr <=  "0011100010110";
		Trees_din <= x"01fe7f20";
		wait for Clk_period;
		Addr <=  "0011100010111";
		Trees_din <= x"28ff1210";
		wait for Clk_period;
		Addr <=  "0011100011000";
		Trees_din <= x"faff7c08";
		wait for Clk_period;
		Addr <=  "0011100011001";
		Trees_din <= x"b0fef104";
		wait for Clk_period;
		Addr <=  "0011100011010";
		Trees_din <= x"ff921d39";
		wait for Clk_period;
		Addr <=  "0011100011011";
		Trees_din <= x"00381d39";
		wait for Clk_period;
		Addr <=  "0011100011100";
		Trees_din <= x"7fff0b04";
		wait for Clk_period;
		Addr <=  "0011100011101";
		Trees_din <= x"00171d39";
		wait for Clk_period;
		Addr <=  "0011100011110";
		Trees_din <= x"ff921d39";
		wait for Clk_period;
		Addr <=  "0011100011111";
		Trees_din <= x"3effc108";
		wait for Clk_period;
		Addr <=  "0011100100000";
		Trees_din <= x"9d004204";
		wait for Clk_period;
		Addr <=  "0011100100001";
		Trees_din <= x"004f1d39";
		wait for Clk_period;
		Addr <=  "0011100100010";
		Trees_din <= x"ffd21d39";
		wait for Clk_period;
		Addr <=  "0011100100011";
		Trees_din <= x"1301d304";
		wait for Clk_period;
		Addr <=  "0011100100100";
		Trees_din <= x"ff8f1d39";
		wait for Clk_period;
		Addr <=  "0011100100101";
		Trees_din <= x"00671d39";
		wait for Clk_period;
		Addr <=  "0011100100110";
		Trees_din <= x"fbff8610";
		wait for Clk_period;
		Addr <=  "0011100100111";
		Trees_din <= x"2bffdf08";
		wait for Clk_period;
		Addr <=  "0011100101000";
		Trees_din <= x"c5ff0c04";
		wait for Clk_period;
		Addr <=  "0011100101001";
		Trees_din <= x"006c1d39";
		wait for Clk_period;
		Addr <=  "0011100101010";
		Trees_din <= x"ffda1d39";
		wait for Clk_period;
		Addr <=  "0011100101011";
		Trees_din <= x"63ff7a04";
		wait for Clk_period;
		Addr <=  "0011100101100";
		Trees_din <= x"ffee1d39";
		wait for Clk_period;
		Addr <=  "0011100101101";
		Trees_din <= x"007a1d39";
		wait for Clk_period;
		Addr <=  "0011100101110";
		Trees_din <= x"59ffdf08";
		wait for Clk_period;
		Addr <=  "0011100101111";
		Trees_din <= x"55002d04";
		wait for Clk_period;
		Addr <=  "0011100110000";
		Trees_din <= x"ffe01d39";
		wait for Clk_period;
		Addr <=  "0011100110001";
		Trees_din <= x"00281d39";
		wait for Clk_period;
		Addr <=  "0011100110010";
		Trees_din <= x"80ffea04";
		wait for Clk_period;
		Addr <=  "0011100110011";
		Trees_din <= x"ff911d39";
		wait for Clk_period;
		Addr <=  "0011100110100";
		Trees_din <= x"003d1d39";
		wait for Clk_period;
		Addr <=  "0011100110101";
		Trees_din <= x"db009418";
		wait for Clk_period;
		Addr <=  "0011100110110";
		Trees_din <= x"dc007a0c";
		wait for Clk_period;
		Addr <=  "0011100110111";
		Trees_din <= x"4400b408";
		wait for Clk_period;
		Addr <=  "0011100111000";
		Trees_din <= x"0a00e004";
		wait for Clk_period;
		Addr <=  "0011100111001";
		Trees_din <= x"ff6a1d39";
		wait for Clk_period;
		Addr <=  "0011100111010";
		Trees_din <= x"ffe01d39";
		wait for Clk_period;
		Addr <=  "0011100111011";
		Trees_din <= x"00161d39";
		wait for Clk_period;
		Addr <=  "0011100111100";
		Trees_din <= x"2bff5f08";
		wait for Clk_period;
		Addr <=  "0011100111101";
		Trees_din <= x"b8ff7604";
		wait for Clk_period;
		Addr <=  "0011100111110";
		Trees_din <= x"000c1d39";
		wait for Clk_period;
		Addr <=  "0011100111111";
		Trees_din <= x"00891d39";
		wait for Clk_period;
		Addr <=  "0011101000000";
		Trees_din <= x"ff9f1d39";
		wait for Clk_period;
		Addr <=  "0011101000001";
		Trees_din <= x"38ffbb14";
		wait for Clk_period;
		Addr <=  "0011101000010";
		Trees_din <= x"15ffa508";
		wait for Clk_period;
		Addr <=  "0011101000011";
		Trees_din <= x"8effb804";
		wait for Clk_period;
		Addr <=  "0011101000100";
		Trees_din <= x"005c1d39";
		wait for Clk_period;
		Addr <=  "0011101000101";
		Trees_din <= x"ff8e1d39";
		wait for Clk_period;
		Addr <=  "0011101000110";
		Trees_din <= x"74ffb904";
		wait for Clk_period;
		Addr <=  "0011101000111";
		Trees_din <= x"ffdf1d39";
		wait for Clk_period;
		Addr <=  "0011101001000";
		Trees_din <= x"b2fffc04";
		wait for Clk_period;
		Addr <=  "0011101001001";
		Trees_din <= x"00b51d39";
		wait for Clk_period;
		Addr <=  "0011101001010";
		Trees_din <= x"00151d39";
		wait for Clk_period;
		Addr <=  "0011101001011";
		Trees_din <= x"83ff7604";
		wait for Clk_period;
		Addr <=  "0011101001100";
		Trees_din <= x"ff8b1d39";
		wait for Clk_period;
		Addr <=  "0011101001101";
		Trees_din <= x"000a1d39";
		wait for Clk_period;
		Addr <=  "0011101001110";
		Trees_din <= x"eaff4348";
		wait for Clk_period;
		Addr <=  "0011101001111";
		Trees_din <= x"40ffeb20";
		wait for Clk_period;
		Addr <=  "0011101010000";
		Trees_din <= x"49003010";
		wait for Clk_period;
		Addr <=  "0011101010001";
		Trees_din <= x"edff3c08";
		wait for Clk_period;
		Addr <=  "0011101010010";
		Trees_din <= x"e2fea904";
		wait for Clk_period;
		Addr <=  "0011101010011";
		Trees_din <= x"00731e75";
		wait for Clk_period;
		Addr <=  "0011101010100";
		Trees_din <= x"ffe51e75";
		wait for Clk_period;
		Addr <=  "0011101010101";
		Trees_din <= x"c800cb04";
		wait for Clk_period;
		Addr <=  "0011101010110";
		Trees_din <= x"ff651e75";
		wait for Clk_period;
		Addr <=  "0011101010111";
		Trees_din <= x"00261e75";
		wait for Clk_period;
		Addr <=  "0011101011000";
		Trees_din <= x"9cffab08";
		wait for Clk_period;
		Addr <=  "0011101011001";
		Trees_din <= x"9affa004";
		wait for Clk_period;
		Addr <=  "0011101011010";
		Trees_din <= x"00001e75";
		wait for Clk_period;
		Addr <=  "0011101011011";
		Trees_din <= x"ff871e75";
		wait for Clk_period;
		Addr <=  "0011101011100";
		Trees_din <= x"fdff2c04";
		wait for Clk_period;
		Addr <=  "0011101011101";
		Trees_din <= x"00931e75";
		wait for Clk_period;
		Addr <=  "0011101011110";
		Trees_din <= x"ffdb1e75";
		wait for Clk_period;
		Addr <=  "0011101011111";
		Trees_din <= x"31ff4708";
		wait for Clk_period;
		Addr <=  "0011101100000";
		Trees_din <= x"09001904";
		wait for Clk_period;
		Addr <=  "0011101100001";
		Trees_din <= x"ff741e75";
		wait for Clk_period;
		Addr <=  "0011101100010";
		Trees_din <= x"002a1e75";
		wait for Clk_period;
		Addr <=  "0011101100011";
		Trees_din <= x"7efee010";
		wait for Clk_period;
		Addr <=  "0011101100100";
		Trees_din <= x"efff8c08";
		wait for Clk_period;
		Addr <=  "0011101100101";
		Trees_din <= x"30001704";
		wait for Clk_period;
		Addr <=  "0011101100110";
		Trees_din <= x"ff871e75";
		wait for Clk_period;
		Addr <=  "0011101100111";
		Trees_din <= x"00221e75";
		wait for Clk_period;
		Addr <=  "0011101101000";
		Trees_din <= x"d2feb204";
		wait for Clk_period;
		Addr <=  "0011101101001";
		Trees_din <= x"ffd31e75";
		wait for Clk_period;
		Addr <=  "0011101101010";
		Trees_din <= x"004f1e75";
		wait for Clk_period;
		Addr <=  "0011101101011";
		Trees_din <= x"93ff8d08";
		wait for Clk_period;
		Addr <=  "0011101101100";
		Trees_din <= x"23ffd004";
		wait for Clk_period;
		Addr <=  "0011101101101";
		Trees_din <= x"ffa91e75";
		wait for Clk_period;
		Addr <=  "0011101101110";
		Trees_din <= x"00661e75";
		wait for Clk_period;
		Addr <=  "0011101101111";
		Trees_din <= x"bfffb704";
		wait for Clk_period;
		Addr <=  "0011101110000";
		Trees_din <= x"00a21e75";
		wait for Clk_period;
		Addr <=  "0011101110001";
		Trees_din <= x"ffa81e75";
		wait for Clk_period;
		Addr <=  "0011101110010";
		Trees_din <= x"c4004040";
		wait for Clk_period;
		Addr <=  "0011101110011";
		Trees_din <= x"6bfe8f20";
		wait for Clk_period;
		Addr <=  "0011101110100";
		Trees_din <= x"64ff0b10";
		wait for Clk_period;
		Addr <=  "0011101110101";
		Trees_din <= x"a6ff8108";
		wait for Clk_period;
		Addr <=  "0011101110110";
		Trees_din <= x"7cff3804";
		wait for Clk_period;
		Addr <=  "0011101110111";
		Trees_din <= x"ffc31e75";
		wait for Clk_period;
		Addr <=  "0011101111000";
		Trees_din <= x"00551e75";
		wait for Clk_period;
		Addr <=  "0011101111001";
		Trees_din <= x"86ff8a04";
		wait for Clk_period;
		Addr <=  "0011101111010";
		Trees_din <= x"ff821e75";
		wait for Clk_period;
		Addr <=  "0011101111011";
		Trees_din <= x"002b1e75";
		wait for Clk_period;
		Addr <=  "0011101111100";
		Trees_din <= x"0dff4208";
		wait for Clk_period;
		Addr <=  "0011101111101";
		Trees_din <= x"39ffd404";
		wait for Clk_period;
		Addr <=  "0011101111110";
		Trees_din <= x"002e1e75";
		wait for Clk_period;
		Addr <=  "0011101111111";
		Trees_din <= x"ffa31e75";
		wait for Clk_period;
		Addr <=  "0011110000000";
		Trees_din <= x"bbffde04";
		wait for Clk_period;
		Addr <=  "0011110000001";
		Trees_din <= x"ff7a1e75";
		wait for Clk_period;
		Addr <=  "0011110000010";
		Trees_din <= x"00541e75";
		wait for Clk_period;
		Addr <=  "0011110000011";
		Trees_din <= x"d9ffd810";
		wait for Clk_period;
		Addr <=  "0011110000100";
		Trees_din <= x"d5ffe608";
		wait for Clk_period;
		Addr <=  "0011110000101";
		Trees_din <= x"1dff9204";
		wait for Clk_period;
		Addr <=  "0011110000110";
		Trees_din <= x"ffbe1e75";
		wait for Clk_period;
		Addr <=  "0011110000111";
		Trees_din <= x"005a1e75";
		wait for Clk_period;
		Addr <=  "0011110001000";
		Trees_din <= x"c3007004";
		wait for Clk_period;
		Addr <=  "0011110001001";
		Trees_din <= x"000c1e75";
		wait for Clk_period;
		Addr <=  "0011110001010";
		Trees_din <= x"00ab1e75";
		wait for Clk_period;
		Addr <=  "0011110001011";
		Trees_din <= x"32fed908";
		wait for Clk_period;
		Addr <=  "0011110001100";
		Trees_din <= x"27001c04";
		wait for Clk_period;
		Addr <=  "0011110001101";
		Trees_din <= x"007f1e75";
		wait for Clk_period;
		Addr <=  "0011110001110";
		Trees_din <= x"ffee1e75";
		wait for Clk_period;
		Addr <=  "0011110001111";
		Trees_din <= x"e5fef104";
		wait for Clk_period;
		Addr <=  "0011110010000";
		Trees_din <= x"003f1e75";
		wait for Clk_period;
		Addr <=  "0011110010001";
		Trees_din <= x"ffd71e75";
		wait for Clk_period;
		Addr <=  "0011110010010";
		Trees_din <= x"9affea14";
		wait for Clk_period;
		Addr <=  "0011110010011";
		Trees_din <= x"e9fef108";
		wait for Clk_period;
		Addr <=  "0011110010100";
		Trees_din <= x"ceffb404";
		wait for Clk_period;
		Addr <=  "0011110010101";
		Trees_din <= x"00571e75";
		wait for Clk_period;
		Addr <=  "0011110010110";
		Trees_din <= x"ff971e75";
		wait for Clk_period;
		Addr <=  "0011110010111";
		Trees_din <= x"dfff0b04";
		wait for Clk_period;
		Addr <=  "0011110011000";
		Trees_din <= x"fffd1e75";
		wait for Clk_period;
		Addr <=  "0011110011001";
		Trees_din <= x"beffbd04";
		wait for Clk_period;
		Addr <=  "0011110011010";
		Trees_din <= x"00251e75";
		wait for Clk_period;
		Addr <=  "0011110011011";
		Trees_din <= x"00d91e75";
		wait for Clk_period;
		Addr <=  "0011110011100";
		Trees_din <= x"ff931e75";
		wait for Clk_period;
		Addr <=  "0011110011101";
		Trees_din <= x"69feb948";
		wait for Clk_period;
		Addr <=  "0011110011110";
		Trees_din <= x"55ffeb20";
		wait for Clk_period;
		Addr <=  "0011110011111";
		Trees_din <= x"cc004518";
		wait for Clk_period;
		Addr <=  "0011110100000";
		Trees_din <= x"10003808";
		wait for Clk_period;
		Addr <=  "0011110100001";
		Trees_din <= x"8800b704";
		wait for Clk_period;
		Addr <=  "0011110100010";
		Trees_din <= x"ff751ff9";
		wait for Clk_period;
		Addr <=  "0011110100011";
		Trees_din <= x"fff01ff9";
		wait for Clk_period;
		Addr <=  "0011110100100";
		Trees_din <= x"d5003d08";
		wait for Clk_period;
		Addr <=  "0011110100101";
		Trees_din <= x"81ff6804";
		wait for Clk_period;
		Addr <=  "0011110100110";
		Trees_din <= x"ffd21ff9";
		wait for Clk_period;
		Addr <=  "0011110100111";
		Trees_din <= x"006a1ff9";
		wait for Clk_period;
		Addr <=  "0011110101000";
		Trees_din <= x"62fed804";
		wait for Clk_period;
		Addr <=  "0011110101001";
		Trees_din <= x"fff31ff9";
		wait for Clk_period;
		Addr <=  "0011110101010";
		Trees_din <= x"ff921ff9";
		wait for Clk_period;
		Addr <=  "0011110101011";
		Trees_din <= x"f7ffa104";
		wait for Clk_period;
		Addr <=  "0011110101100";
		Trees_din <= x"00961ff9";
		wait for Clk_period;
		Addr <=  "0011110101101";
		Trees_din <= x"00031ff9";
		wait for Clk_period;
		Addr <=  "0011110101110";
		Trees_din <= x"0800d418";
		wait for Clk_period;
		Addr <=  "0011110101111";
		Trees_din <= x"42fff810";
		wait for Clk_period;
		Addr <=  "0011110110000";
		Trees_din <= x"4cfee208";
		wait for Clk_period;
		Addr <=  "0011110110001";
		Trees_din <= x"8e004004";
		wait for Clk_period;
		Addr <=  "0011110110010";
		Trees_din <= x"ff941ff9";
		wait for Clk_period;
		Addr <=  "0011110110011";
		Trees_din <= x"00621ff9";
		wait for Clk_period;
		Addr <=  "0011110110100";
		Trees_din <= x"77fe7404";
		wait for Clk_period;
		Addr <=  "0011110110101";
		Trees_din <= x"ffd41ff9";
		wait for Clk_period;
		Addr <=  "0011110110110";
		Trees_din <= x"00961ff9";
		wait for Clk_period;
		Addr <=  "0011110110111";
		Trees_din <= x"71fed004";
		wait for Clk_period;
		Addr <=  "0011110111000";
		Trees_din <= x"00311ff9";
		wait for Clk_period;
		Addr <=  "0011110111001";
		Trees_din <= x"ff951ff9";
		wait for Clk_period;
		Addr <=  "0011110111010";
		Trees_din <= x"86000b08";
		wait for Clk_period;
		Addr <=  "0011110111011";
		Trees_din <= x"88008504";
		wait for Clk_period;
		Addr <=  "0011110111100";
		Trees_din <= x"ff891ff9";
		wait for Clk_period;
		Addr <=  "0011110111101";
		Trees_din <= x"00211ff9";
		wait for Clk_period;
		Addr <=  "0011110111110";
		Trees_din <= x"d3fe8c04";
		wait for Clk_period;
		Addr <=  "0011110111111";
		Trees_din <= x"00741ff9";
		wait for Clk_period;
		Addr <=  "0011111000000";
		Trees_din <= x"00181ff9";
		wait for Clk_period;
		Addr <=  "0011111000001";
		Trees_din <= x"99ff1240";
		wait for Clk_period;
		Addr <=  "0011111000010";
		Trees_din <= x"01fec620";
		wait for Clk_period;
		Addr <=  "0011111000011";
		Trees_din <= x"9bff2910";
		wait for Clk_period;
		Addr <=  "0011111000100";
		Trees_din <= x"44000d08";
		wait for Clk_period;
		Addr <=  "0011111000101";
		Trees_din <= x"6effff04";
		wait for Clk_period;
		Addr <=  "0011111000110";
		Trees_din <= x"fffb1ff9";
		wait for Clk_period;
		Addr <=  "0011111000111";
		Trees_din <= x"00611ff9";
		wait for Clk_period;
		Addr <=  "0011111001000";
		Trees_din <= x"67ff3004";
		wait for Clk_period;
		Addr <=  "0011111001001";
		Trees_din <= x"00301ff9";
		wait for Clk_period;
		Addr <=  "0011111001010";
		Trees_din <= x"ffad1ff9";
		wait for Clk_period;
		Addr <=  "0011111001011";
		Trees_din <= x"5a00b308";
		wait for Clk_period;
		Addr <=  "0011111001100";
		Trees_din <= x"29ff4304";
		wait for Clk_period;
		Addr <=  "0011111001101";
		Trees_din <= x"ffbb1ff9";
		wait for Clk_period;
		Addr <=  "0011111001110";
		Trees_din <= x"00161ff9";
		wait for Clk_period;
		Addr <=  "0011111001111";
		Trees_din <= x"e9fe1504";
		wait for Clk_period;
		Addr <=  "0011111010000";
		Trees_din <= x"00271ff9";
		wait for Clk_period;
		Addr <=  "0011111010001";
		Trees_din <= x"ff761ff9";
		wait for Clk_period;
		Addr <=  "0011111010010";
		Trees_din <= x"d2fee110";
		wait for Clk_period;
		Addr <=  "0011111010011";
		Trees_din <= x"9afef408";
		wait for Clk_period;
		Addr <=  "0011111010100";
		Trees_din <= x"f4fea504";
		wait for Clk_period;
		Addr <=  "0011111010101";
		Trees_din <= x"00a01ff9";
		wait for Clk_period;
		Addr <=  "0011111010110";
		Trees_din <= x"ffe81ff9";
		wait for Clk_period;
		Addr <=  "0011111010111";
		Trees_din <= x"2aff1404";
		wait for Clk_period;
		Addr <=  "0011111011000";
		Trees_din <= x"00821ff9";
		wait for Clk_period;
		Addr <=  "0011111011001";
		Trees_din <= x"ff8b1ff9";
		wait for Clk_period;
		Addr <=  "0011111011010";
		Trees_din <= x"50ff9f08";
		wait for Clk_period;
		Addr <=  "0011111011011";
		Trees_din <= x"f1ff7004";
		wait for Clk_period;
		Addr <=  "0011111011100";
		Trees_din <= x"00361ff9";
		wait for Clk_period;
		Addr <=  "0011111011101";
		Trees_din <= x"ff8b1ff9";
		wait for Clk_period;
		Addr <=  "0011111011110";
		Trees_din <= x"c5ff3704";
		wait for Clk_period;
		Addr <=  "0011111011111";
		Trees_din <= x"ffcb1ff9";
		wait for Clk_period;
		Addr <=  "0011111100000";
		Trees_din <= x"00871ff9";
		wait for Clk_period;
		Addr <=  "0011111100001";
		Trees_din <= x"5400341c";
		wait for Clk_period;
		Addr <=  "0011111100010";
		Trees_din <= x"6cffc910";
		wait for Clk_period;
		Addr <=  "0011111100011";
		Trees_din <= x"9a000e08";
		wait for Clk_period;
		Addr <=  "0011111100100";
		Trees_din <= x"06fef204";
		wait for Clk_period;
		Addr <=  "0011111100101";
		Trees_din <= x"ff8d1ff9";
		wait for Clk_period;
		Addr <=  "0011111100110";
		Trees_din <= x"00361ff9";
		wait for Clk_period;
		Addr <=  "0011111100111";
		Trees_din <= x"0b002404";
		wait for Clk_period;
		Addr <=  "0011111101000";
		Trees_din <= x"ff781ff9";
		wait for Clk_period;
		Addr <=  "0011111101001";
		Trees_din <= x"00171ff9";
		wait for Clk_period;
		Addr <=  "0011111101010";
		Trees_din <= x"adfef204";
		wait for Clk_period;
		Addr <=  "0011111101011";
		Trees_din <= x"00201ff9";
		wait for Clk_period;
		Addr <=  "0011111101100";
		Trees_din <= x"31005204";
		wait for Clk_period;
		Addr <=  "0011111101101";
		Trees_din <= x"ff6e1ff9";
		wait for Clk_period;
		Addr <=  "0011111101110";
		Trees_din <= x"ffeb1ff9";
		wait for Clk_period;
		Addr <=  "0011111101111";
		Trees_din <= x"5ffec810";
		wait for Clk_period;
		Addr <=  "0011111110000";
		Trees_din <= x"6afff108";
		wait for Clk_period;
		Addr <=  "0011111110001";
		Trees_din <= x"a9fe4604";
		wait for Clk_period;
		Addr <=  "0011111110010";
		Trees_din <= x"00701ff9";
		wait for Clk_period;
		Addr <=  "0011111110011";
		Trees_din <= x"ff781ff9";
		wait for Clk_period;
		Addr <=  "0011111110100";
		Trees_din <= x"1cff2c04";
		wait for Clk_period;
		Addr <=  "0011111110101";
		Trees_din <= x"009b1ff9";
		wait for Clk_period;
		Addr <=  "0011111110110";
		Trees_din <= x"ffcc1ff9";
		wait for Clk_period;
		Addr <=  "0011111110111";
		Trees_din <= x"2bffc408";
		wait for Clk_period;
		Addr <=  "0011111111000";
		Trees_din <= x"77feda04";
		wait for Clk_period;
		Addr <=  "0011111111001";
		Trees_din <= x"00761ff9";
		wait for Clk_period;
		Addr <=  "0011111111010";
		Trees_din <= x"ffda1ff9";
		wait for Clk_period;
		Addr <=  "0011111111011";
		Trees_din <= x"eaff3c04";
		wait for Clk_period;
		Addr <=  "0011111111100";
		Trees_din <= x"fff01ff9";
		wait for Clk_period;
		Addr <=  "0011111111101";
		Trees_din <= x"00951ff9";
		wait for Clk_period;
		Addr <=  "0011111111110";
		Trees_din <= x"6f003e74";
		wait for Clk_period;
		Addr <=  "0011111111111";
		Trees_din <= x"36ffc838";
		wait for Clk_period;
		Addr <=  "0100000000000";
		Trees_din <= x"00feff18";
		wait for Clk_period;
		Addr <=  "0100000000001";
		Trees_din <= x"c3ff3708";
		wait for Clk_period;
		Addr <=  "0100000000010";
		Trees_din <= x"7aff6104";
		wait for Clk_period;
		Addr <=  "0100000000011";
		Trees_din <= x"00b720f5";
		wait for Clk_period;
		Addr <=  "0100000000100";
		Trees_din <= x"001220f5";
		wait for Clk_period;
		Addr <=  "0100000000101";
		Trees_din <= x"82fe7f08";
		wait for Clk_period;
		Addr <=  "0100000000110";
		Trees_din <= x"21ffe404";
		wait for Clk_period;
		Addr <=  "0100000000111";
		Trees_din <= x"001220f5";
		wait for Clk_period;
		Addr <=  "0100000001000";
		Trees_din <= x"007620f5";
		wait for Clk_period;
		Addr <=  "0100000001001";
		Trees_din <= x"2aff7204";
		wait for Clk_period;
		Addr <=  "0100000001010";
		Trees_din <= x"001820f5";
		wait for Clk_period;
		Addr <=  "0100000001011";
		Trees_din <= x"ff9220f5";
		wait for Clk_period;
		Addr <=  "0100000001100";
		Trees_din <= x"3eff6810";
		wait for Clk_period;
		Addr <=  "0100000001101";
		Trees_din <= x"b4fee908";
		wait for Clk_period;
		Addr <=  "0100000001110";
		Trees_din <= x"d8004804";
		wait for Clk_period;
		Addr <=  "0100000001111";
		Trees_din <= x"003f20f5";
		wait for Clk_period;
		Addr <=  "0100000010000";
		Trees_din <= x"ffef20f5";
		wait for Clk_period;
		Addr <=  "0100000010001";
		Trees_din <= x"4cffa104";
		wait for Clk_period;
		Addr <=  "0100000010010";
		Trees_din <= x"ffd320f5";
		wait for Clk_period;
		Addr <=  "0100000010011";
		Trees_din <= x"003b20f5";
		wait for Clk_period;
		Addr <=  "0100000010100";
		Trees_din <= x"fcfebd08";
		wait for Clk_period;
		Addr <=  "0100000010101";
		Trees_din <= x"11ff6604";
		wait for Clk_period;
		Addr <=  "0100000010110";
		Trees_din <= x"ff7720f5";
		wait for Clk_period;
		Addr <=  "0100000010111";
		Trees_din <= x"000f20f5";
		wait for Clk_period;
		Addr <=  "0100000011000";
		Trees_din <= x"8bffbd04";
		wait for Clk_period;
		Addr <=  "0100000011001";
		Trees_din <= x"ffe220f5";
		wait for Clk_period;
		Addr <=  "0100000011010";
		Trees_din <= x"003b20f5";
		wait for Clk_period;
		Addr <=  "0100000011011";
		Trees_din <= x"0efea620";
		wait for Clk_period;
		Addr <=  "0100000011100";
		Trees_din <= x"c7feee10";
		wait for Clk_period;
		Addr <=  "0100000011101";
		Trees_din <= x"8a001408";
		wait for Clk_period;
		Addr <=  "0100000011110";
		Trees_din <= x"beff5604";
		wait for Clk_period;
		Addr <=  "0100000011111";
		Trees_din <= x"002e20f5";
		wait for Clk_period;
		Addr <=  "0100000100000";
		Trees_din <= x"ff7020f5";
		wait for Clk_period;
		Addr <=  "0100000100001";
		Trees_din <= x"6aff6e04";
		wait for Clk_period;
		Addr <=  "0100000100010";
		Trees_din <= x"009920f5";
		wait for Clk_period;
		Addr <=  "0100000100011";
		Trees_din <= x"ffe320f5";
		wait for Clk_period;
		Addr <=  "0100000100100";
		Trees_din <= x"fcff6108";
		wait for Clk_period;
		Addr <=  "0100000100101";
		Trees_din <= x"a1fea904";
		wait for Clk_period;
		Addr <=  "0100000100110";
		Trees_din <= x"ffbe20f5";
		wait for Clk_period;
		Addr <=  "0100000100111";
		Trees_din <= x"008820f5";
		wait for Clk_period;
		Addr <=  "0100000101000";
		Trees_din <= x"3efef804";
		wait for Clk_period;
		Addr <=  "0100000101001";
		Trees_din <= x"005b20f5";
		wait for Clk_period;
		Addr <=  "0100000101010";
		Trees_din <= x"ff8e20f5";
		wait for Clk_period;
		Addr <=  "0100000101011";
		Trees_din <= x"49ff740c";
		wait for Clk_period;
		Addr <=  "0100000101100";
		Trees_din <= x"96ff4708";
		wait for Clk_period;
		Addr <=  "0100000101101";
		Trees_din <= x"0eff4b04";
		wait for Clk_period;
		Addr <=  "0100000101110";
		Trees_din <= x"fffd20f5";
		wait for Clk_period;
		Addr <=  "0100000101111";
		Trees_din <= x"007f20f5";
		wait for Clk_period;
		Addr <=  "0100000110000";
		Trees_din <= x"ffa220f5";
		wait for Clk_period;
		Addr <=  "0100000110001";
		Trees_din <= x"2cff1208";
		wait for Clk_period;
		Addr <=  "0100000110010";
		Trees_din <= x"d1ff1204";
		wait for Clk_period;
		Addr <=  "0100000110011";
		Trees_din <= x"006d20f5";
		wait for Clk_period;
		Addr <=  "0100000110100";
		Trees_din <= x"ffa820f5";
		wait for Clk_period;
		Addr <=  "0100000110101";
		Trees_din <= x"17ff5e04";
		wait for Clk_period;
		Addr <=  "0100000110110";
		Trees_din <= x"000720f5";
		wait for Clk_period;
		Addr <=  "0100000110111";
		Trees_din <= x"ff6820f5";
		wait for Clk_period;
		Addr <=  "0100000111000";
		Trees_din <= x"3eff1a04";
		wait for Clk_period;
		Addr <=  "0100000111001";
		Trees_din <= x"003d20f5";
		wait for Clk_period;
		Addr <=  "0100000111010";
		Trees_din <= x"c1ff8704";
		wait for Clk_period;
		Addr <=  "0100000111011";
		Trees_din <= x"ff7220f5";
		wait for Clk_period;
		Addr <=  "0100000111100";
		Trees_din <= x"000a20f5";
		wait for Clk_period;
		Addr <=  "0100000111101";
		Trees_din <= x"a4ff1b38";
		wait for Clk_period;
		Addr <=  "0100000111110";
		Trees_din <= x"fcfec508";
		wait for Clk_period;
		Addr <=  "0100000111111";
		Trees_din <= x"a5ff6704";
		wait for Clk_period;
		Addr <=  "0100001000000";
		Trees_din <= x"ff8d2249";
		wait for Clk_period;
		Addr <=  "0100001000001";
		Trees_din <= x"fff32249";
		wait for Clk_period;
		Addr <=  "0100001000010";
		Trees_din <= x"95ff2718";
		wait for Clk_period;
		Addr <=  "0100001000011";
		Trees_din <= x"88ffce08";
		wait for Clk_period;
		Addr <=  "0100001000100";
		Trees_din <= x"8affc404";
		wait for Clk_period;
		Addr <=  "0100001000101";
		Trees_din <= x"ff7c2249";
		wait for Clk_period;
		Addr <=  "0100001000110";
		Trees_din <= x"001a2249";
		wait for Clk_period;
		Addr <=  "0100001000111";
		Trees_din <= x"f9ff4408";
		wait for Clk_period;
		Addr <=  "0100001001000";
		Trees_din <= x"14fed604";
		wait for Clk_period;
		Addr <=  "0100001001001";
		Trees_din <= x"ffe62249";
		wait for Clk_period;
		Addr <=  "0100001001010";
		Trees_din <= x"00852249";
		wait for Clk_period;
		Addr <=  "0100001001011";
		Trees_din <= x"a6ff1104";
		wait for Clk_period;
		Addr <=  "0100001001100";
		Trees_din <= x"004b2249";
		wait for Clk_period;
		Addr <=  "0100001001101";
		Trees_din <= x"ff882249";
		wait for Clk_period;
		Addr <=  "0100001001110";
		Trees_din <= x"1eff900c";
		wait for Clk_period;
		Addr <=  "0100001001111";
		Trees_din <= x"f2024c04";
		wait for Clk_period;
		Addr <=  "0100001010000";
		Trees_din <= x"ff902249";
		wait for Clk_period;
		Addr <=  "0100001010001";
		Trees_din <= x"b8ff7904";
		wait for Clk_period;
		Addr <=  "0100001010010";
		Trees_din <= x"006d2249";
		wait for Clk_period;
		Addr <=  "0100001010011";
		Trees_din <= x"ffce2249";
		wait for Clk_period;
		Addr <=  "0100001010100";
		Trees_din <= x"fdff0a04";
		wait for Clk_period;
		Addr <=  "0100001010101";
		Trees_din <= x"ffc12249";
		wait for Clk_period;
		Addr <=  "0100001010110";
		Trees_din <= x"cbffa504";
		wait for Clk_period;
		Addr <=  "0100001010111";
		Trees_din <= x"002b2249";
		wait for Clk_period;
		Addr <=  "0100001011000";
		Trees_din <= x"00d32249";
		wait for Clk_period;
		Addr <=  "0100001011001";
		Trees_din <= x"21ffb33c";
		wait for Clk_period;
		Addr <=  "0100001011010";
		Trees_din <= x"14ff2e20";
		wait for Clk_period;
		Addr <=  "0100001011011";
		Trees_din <= x"3aff3d10";
		wait for Clk_period;
		Addr <=  "0100001011100";
		Trees_din <= x"a9fff808";
		wait for Clk_period;
		Addr <=  "0100001011101";
		Trees_din <= x"61fee704";
		wait for Clk_period;
		Addr <=  "0100001011110";
		Trees_din <= x"fff82249";
		wait for Clk_period;
		Addr <=  "0100001011111";
		Trees_din <= x"00562249";
		wait for Clk_period;
		Addr <=  "0100001100000";
		Trees_din <= x"45ff3204";
		wait for Clk_period;
		Addr <=  "0100001100001";
		Trees_din <= x"ff912249";
		wait for Clk_period;
		Addr <=  "0100001100010";
		Trees_din <= x"002e2249";
		wait for Clk_period;
		Addr <=  "0100001100011";
		Trees_din <= x"05003708";
		wait for Clk_period;
		Addr <=  "0100001100100";
		Trees_din <= x"20ff8204";
		wait for Clk_period;
		Addr <=  "0100001100101";
		Trees_din <= x"ffbd2249";
		wait for Clk_period;
		Addr <=  "0100001100110";
		Trees_din <= x"005e2249";
		wait for Clk_period;
		Addr <=  "0100001100111";
		Trees_din <= x"69fef504";
		wait for Clk_period;
		Addr <=  "0100001101000";
		Trees_din <= x"00212249";
		wait for Clk_period;
		Addr <=  "0100001101001";
		Trees_din <= x"ffa82249";
		wait for Clk_period;
		Addr <=  "0100001101010";
		Trees_din <= x"9affe710";
		wait for Clk_period;
		Addr <=  "0100001101011";
		Trees_din <= x"34ffef08";
		wait for Clk_period;
		Addr <=  "0100001101100";
		Trees_din <= x"b3fedf04";
		wait for Clk_period;
		Addr <=  "0100001101101";
		Trees_din <= x"ffb22249";
		wait for Clk_period;
		Addr <=  "0100001101110";
		Trees_din <= x"005d2249";
		wait for Clk_period;
		Addr <=  "0100001101111";
		Trees_din <= x"7efe7404";
		wait for Clk_period;
		Addr <=  "0100001110000";
		Trees_din <= x"001c2249";
		wait for Clk_period;
		Addr <=  "0100001110001";
		Trees_din <= x"ff9e2249";
		wait for Clk_period;
		Addr <=  "0100001110010";
		Trees_din <= x"c7001d08";
		wait for Clk_period;
		Addr <=  "0100001110011";
		Trees_din <= x"aa001b04";
		wait for Clk_period;
		Addr <=  "0100001110100";
		Trees_din <= x"ff742249";
		wait for Clk_period;
		Addr <=  "0100001110101";
		Trees_din <= x"00112249";
		wait for Clk_period;
		Addr <=  "0100001110110";
		Trees_din <= x"006c2249";
		wait for Clk_period;
		Addr <=  "0100001110111";
		Trees_din <= x"12ff571c";
		wait for Clk_period;
		Addr <=  "0100001111000";
		Trees_din <= x"ab00940c";
		wait for Clk_period;
		Addr <=  "0100001111001";
		Trees_din <= x"1f00c408";
		wait for Clk_period;
		Addr <=  "0100001111010";
		Trees_din <= x"64fe6704";
		wait for Clk_period;
		Addr <=  "0100001111011";
		Trees_din <= x"fff42249";
		wait for Clk_period;
		Addr <=  "0100001111100";
		Trees_din <= x"ff692249";
		wait for Clk_period;
		Addr <=  "0100001111101";
		Trees_din <= x"000c2249";
		wait for Clk_period;
		Addr <=  "0100001111110";
		Trees_din <= x"7ffef608";
		wait for Clk_period;
		Addr <=  "0100001111111";
		Trees_din <= x"06003304";
		wait for Clk_period;
		Addr <=  "0100010000000";
		Trees_din <= x"00952249";
		wait for Clk_period;
		Addr <=  "0100010000001";
		Trees_din <= x"ffd32249";
		wait for Clk_period;
		Addr <=  "0100010000010";
		Trees_din <= x"98fe4404";
		wait for Clk_period;
		Addr <=  "0100010000011";
		Trees_din <= x"003f2249";
		wait for Clk_period;
		Addr <=  "0100010000100";
		Trees_din <= x"ff7b2249";
		wait for Clk_period;
		Addr <=  "0100010000101";
		Trees_din <= x"15fee60c";
		wait for Clk_period;
		Addr <=  "0100010000110";
		Trees_din <= x"79ff0d04";
		wait for Clk_period;
		Addr <=  "0100010000111";
		Trees_din <= x"ffa12249";
		wait for Clk_period;
		Addr <=  "0100010001000";
		Trees_din <= x"eeffdf04";
		wait for Clk_period;
		Addr <=  "0100010001001";
		Trees_din <= x"fff62249";
		wait for Clk_period;
		Addr <=  "0100010001010";
		Trees_din <= x"00cc2249";
		wait for Clk_period;
		Addr <=  "0100010001011";
		Trees_din <= x"33fef408";
		wait for Clk_period;
		Addr <=  "0100010001100";
		Trees_din <= x"af001104";
		wait for Clk_period;
		Addr <=  "0100010001101";
		Trees_din <= x"ffa02249";
		wait for Clk_period;
		Addr <=  "0100010001110";
		Trees_din <= x"00162249";
		wait for Clk_period;
		Addr <=  "0100010001111";
		Trees_din <= x"33ffc804";
		wait for Clk_period;
		Addr <=  "0100010010000";
		Trees_din <= x"00102249";
		wait for Clk_period;
		Addr <=  "0100010010001";
		Trees_din <= x"ffaa2249";
		wait for Clk_period;
		Addr <=  "0100010010010";
		Trees_din <= x"1f011f6c";
		wait for Clk_period;
		Addr <=  "0100010010011";
		Trees_din <= x"99ff1340";
		wait for Clk_period;
		Addr <=  "0100010010100";
		Trees_din <= x"d9ffc620";
		wait for Clk_period;
		Addr <=  "0100010010101";
		Trees_din <= x"93ff9f10";
		wait for Clk_period;
		Addr <=  "0100010010110";
		Trees_din <= x"f0ffbb08";
		wait for Clk_period;
		Addr <=  "0100010010111";
		Trees_din <= x"9c002604";
		wait for Clk_period;
		Addr <=  "0100010011000";
		Trees_din <= x"ff992355";
		wait for Clk_period;
		Addr <=  "0100010011001";
		Trees_din <= x"003d2355";
		wait for Clk_period;
		Addr <=  "0100010011010";
		Trees_din <= x"37ff5c04";
		wait for Clk_period;
		Addr <=  "0100010011011";
		Trees_din <= x"00572355";
		wait for Clk_period;
		Addr <=  "0100010011100";
		Trees_din <= x"ffae2355";
		wait for Clk_period;
		Addr <=  "0100010011101";
		Trees_din <= x"f9ff5908";
		wait for Clk_period;
		Addr <=  "0100010011110";
		Trees_din <= x"46fee504";
		wait for Clk_period;
		Addr <=  "0100010011111";
		Trees_din <= x"000e2355";
		wait for Clk_period;
		Addr <=  "0100010100000";
		Trees_din <= x"ffa02355";
		wait for Clk_period;
		Addr <=  "0100010100001";
		Trees_din <= x"e9febe04";
		wait for Clk_period;
		Addr <=  "0100010100010";
		Trees_din <= x"ffc62355";
		wait for Clk_period;
		Addr <=  "0100010100011";
		Trees_din <= x"00672355";
		wait for Clk_period;
		Addr <=  "0100010100100";
		Trees_din <= x"77fef310";
		wait for Clk_period;
		Addr <=  "0100010100101";
		Trees_din <= x"5a007908";
		wait for Clk_period;
		Addr <=  "0100010100110";
		Trees_din <= x"5cffea04";
		wait for Clk_period;
		Addr <=  "0100010100111";
		Trees_din <= x"00482355";
		wait for Clk_period;
		Addr <=  "0100010101000";
		Trees_din <= x"ffd22355";
		wait for Clk_period;
		Addr <=  "0100010101001";
		Trees_din <= x"f4fe3504";
		wait for Clk_period;
		Addr <=  "0100010101010";
		Trees_din <= x"00422355";
		wait for Clk_period;
		Addr <=  "0100010101011";
		Trees_din <= x"ff842355";
		wait for Clk_period;
		Addr <=  "0100010101100";
		Trees_din <= x"e5ff3d08";
		wait for Clk_period;
		Addr <=  "0100010101101";
		Trees_din <= x"0400cf04";
		wait for Clk_period;
		Addr <=  "0100010101110";
		Trees_din <= x"00402355";
		wait for Clk_period;
		Addr <=  "0100010101111";
		Trees_din <= x"ffca2355";
		wait for Clk_period;
		Addr <=  "0100010110000";
		Trees_din <= x"42ff3904";
		wait for Clk_period;
		Addr <=  "0100010110001";
		Trees_din <= x"00292355";
		wait for Clk_period;
		Addr <=  "0100010110010";
		Trees_din <= x"ff7b2355";
		wait for Clk_period;
		Addr <=  "0100010110011";
		Trees_din <= x"f9fe7510";
		wait for Clk_period;
		Addr <=  "0100010110100";
		Trees_din <= x"01fe1c08";
		wait for Clk_period;
		Addr <=  "0100010110101";
		Trees_din <= x"b5ff1b04";
		wait for Clk_period;
		Addr <=  "0100010110110";
		Trees_din <= x"ffe72355";
		wait for Clk_period;
		Addr <=  "0100010110111";
		Trees_din <= x"00552355";
		wait for Clk_period;
		Addr <=  "0100010111000";
		Trees_din <= x"92ff8e04";
		wait for Clk_period;
		Addr <=  "0100010111001";
		Trees_din <= x"ff712355";
		wait for Clk_period;
		Addr <=  "0100010111010";
		Trees_din <= x"fff52355";
		wait for Clk_period;
		Addr <=  "0100010111011";
		Trees_din <= x"c6ffe610";
		wait for Clk_period;
		Addr <=  "0100010111100";
		Trees_din <= x"36ffa208";
		wait for Clk_period;
		Addr <=  "0100010111101";
		Trees_din <= x"49000704";
		wait for Clk_period;
		Addr <=  "0100010111110";
		Trees_din <= x"004b2355";
		wait for Clk_period;
		Addr <=  "0100010111111";
		Trees_din <= x"00022355";
		wait for Clk_period;
		Addr <=  "0100011000000";
		Trees_din <= x"5dffe104";
		wait for Clk_period;
		Addr <=  "0100011000001";
		Trees_din <= x"ffb22355";
		wait for Clk_period;
		Addr <=  "0100011000010";
		Trees_din <= x"00272355";
		wait for Clk_period;
		Addr <=  "0100011000011";
		Trees_din <= x"ce003608";
		wait for Clk_period;
		Addr <=  "0100011000100";
		Trees_din <= x"69fed204";
		wait for Clk_period;
		Addr <=  "0100011000101";
		Trees_din <= x"fffd2355";
		wait for Clk_period;
		Addr <=  "0100011000110";
		Trees_din <= x"ff762355";
		wait for Clk_period;
		Addr <=  "0100011000111";
		Trees_din <= x"00482355";
		wait for Clk_period;
		Addr <=  "0100011001000";
		Trees_din <= x"bdffca10";
		wait for Clk_period;
		Addr <=  "0100011001001";
		Trees_din <= x"d600fe0c";
		wait for Clk_period;
		Addr <=  "0100011001010";
		Trees_din <= x"66ff9508";
		wait for Clk_period;
		Addr <=  "0100011001011";
		Trees_din <= x"70fecb04";
		wait for Clk_period;
		Addr <=  "0100011001100";
		Trees_din <= x"ffae2355";
		wait for Clk_period;
		Addr <=  "0100011001101";
		Trees_din <= x"00462355";
		wait for Clk_period;
		Addr <=  "0100011001110";
		Trees_din <= x"00922355";
		wait for Clk_period;
		Addr <=  "0100011001111";
		Trees_din <= x"ffd62355";
		wait for Clk_period;
		Addr <=  "0100011010000";
		Trees_din <= x"a2ffca04";
		wait for Clk_period;
		Addr <=  "0100011010001";
		Trees_din <= x"ff892355";
		wait for Clk_period;
		Addr <=  "0100011010010";
		Trees_din <= x"8ffeff04";
		wait for Clk_period;
		Addr <=  "0100011010011";
		Trees_din <= x"00632355";
		wait for Clk_period;
		Addr <=  "0100011010100";
		Trees_din <= x"ffef2355";
		wait for Clk_period;
		Addr <=  "0100011010101";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0100011010110";
		Trees_din <= x"43ffe068";
		wait for Clk_period;
		Addr <=  "0100011010111";
		Trees_din <= x"19ffa03c";
		wait for Clk_period;
		Addr <=  "0100011011000";
		Trees_din <= x"9dff511c";
		wait for Clk_period;
		Addr <=  "0100011011001";
		Trees_din <= x"28fec00c";
		wait for Clk_period;
		Addr <=  "0100011011010";
		Trees_din <= x"87ffca08";
		wait for Clk_period;
		Addr <=  "0100011011011";
		Trees_din <= x"89009e04";
		wait for Clk_period;
		Addr <=  "0100011011100";
		Trees_din <= x"ff702495";
		wait for Clk_period;
		Addr <=  "0100011011101";
		Trees_din <= x"ffef2495";
		wait for Clk_period;
		Addr <=  "0100011011110";
		Trees_din <= x"003a2495";
		wait for Clk_period;
		Addr <=  "0100011011111";
		Trees_din <= x"cafed708";
		wait for Clk_period;
		Addr <=  "0100011100000";
		Trees_din <= x"69fed804";
		wait for Clk_period;
		Addr <=  "0100011100001";
		Trees_din <= x"00562495";
		wait for Clk_period;
		Addr <=  "0100011100010";
		Trees_din <= x"fff72495";
		wait for Clk_period;
		Addr <=  "0100011100011";
		Trees_din <= x"57ff7a04";
		wait for Clk_period;
		Addr <=  "0100011100100";
		Trees_din <= x"ff782495";
		wait for Clk_period;
		Addr <=  "0100011100101";
		Trees_din <= x"00282495";
		wait for Clk_period;
		Addr <=  "0100011100110";
		Trees_din <= x"d3ff7610";
		wait for Clk_period;
		Addr <=  "0100011100111";
		Trees_din <= x"6d001808";
		wait for Clk_period;
		Addr <=  "0100011101000";
		Trees_din <= x"90ff6504";
		wait for Clk_period;
		Addr <=  "0100011101001";
		Trees_din <= x"ffcc2495";
		wait for Clk_period;
		Addr <=  "0100011101010";
		Trees_din <= x"00232495";
		wait for Clk_period;
		Addr <=  "0100011101011";
		Trees_din <= x"70ff1404";
		wait for Clk_period;
		Addr <=  "0100011101100";
		Trees_din <= x"00172495";
		wait for Clk_period;
		Addr <=  "0100011101101";
		Trees_din <= x"00592495";
		wait for Clk_period;
		Addr <=  "0100011101110";
		Trees_din <= x"2bff3208";
		wait for Clk_period;
		Addr <=  "0100011101111";
		Trees_din <= x"ceff9104";
		wait for Clk_period;
		Addr <=  "0100011110000";
		Trees_din <= x"00722495";
		wait for Clk_period;
		Addr <=  "0100011110001";
		Trees_din <= x"ffb02495";
		wait for Clk_period;
		Addr <=  "0100011110010";
		Trees_din <= x"a2ff3304";
		wait for Clk_period;
		Addr <=  "0100011110011";
		Trees_din <= x"003b2495";
		wait for Clk_period;
		Addr <=  "0100011110100";
		Trees_din <= x"ff862495";
		wait for Clk_period;
		Addr <=  "0100011110101";
		Trees_din <= x"db00ac18";
		wait for Clk_period;
		Addr <=  "0100011110110";
		Trees_din <= x"35fe8510";
		wait for Clk_period;
		Addr <=  "0100011110111";
		Trees_din <= x"28fee708";
		wait for Clk_period;
		Addr <=  "0100011111000";
		Trees_din <= x"4bff0104";
		wait for Clk_period;
		Addr <=  "0100011111001";
		Trees_din <= x"00102495";
		wait for Clk_period;
		Addr <=  "0100011111010";
		Trees_din <= x"00682495";
		wait for Clk_period;
		Addr <=  "0100011111011";
		Trees_din <= x"11ff8204";
		wait for Clk_period;
		Addr <=  "0100011111100";
		Trees_din <= x"ff9a2495";
		wait for Clk_period;
		Addr <=  "0100011111101";
		Trees_din <= x"00012495";
		wait for Clk_period;
		Addr <=  "0100011111110";
		Trees_din <= x"51007704";
		wait for Clk_period;
		Addr <=  "0100011111111";
		Trees_din <= x"ff712495";
		wait for Clk_period;
		Addr <=  "0100100000000";
		Trees_din <= x"ffea2495";
		wait for Clk_period;
		Addr <=  "0100100000001";
		Trees_din <= x"aaff7810";
		wait for Clk_period;
		Addr <=  "0100100000010";
		Trees_din <= x"f1ff9c08";
		wait for Clk_period;
		Addr <=  "0100100000011";
		Trees_din <= x"71ff0d04";
		wait for Clk_period;
		Addr <=  "0100100000100";
		Trees_din <= x"008a2495";
		wait for Clk_period;
		Addr <=  "0100100000101";
		Trees_din <= x"002a2495";
		wait for Clk_period;
		Addr <=  "0100100000110";
		Trees_din <= x"20005604";
		wait for Clk_period;
		Addr <=  "0100100000111";
		Trees_din <= x"ffb02495";
		wait for Clk_period;
		Addr <=  "0100100001000";
		Trees_din <= x"00302495";
		wait for Clk_period;
		Addr <=  "0100100001001";
		Trees_din <= x"ffa92495";
		wait for Clk_period;
		Addr <=  "0100100001010";
		Trees_din <= x"a9feae0c";
		wait for Clk_period;
		Addr <=  "0100100001011";
		Trees_din <= x"a4ff1404";
		wait for Clk_period;
		Addr <=  "0100100001100";
		Trees_din <= x"00b02495";
		wait for Clk_period;
		Addr <=  "0100100001101";
		Trees_din <= x"8ffeea04";
		wait for Clk_period;
		Addr <=  "0100100001110";
		Trees_din <= x"00402495";
		wait for Clk_period;
		Addr <=  "0100100001111";
		Trees_din <= x"ffa72495";
		wait for Clk_period;
		Addr <=  "0100100010000";
		Trees_din <= x"75005c14";
		wait for Clk_period;
		Addr <=  "0100100010001";
		Trees_din <= x"5e007a10";
		wait for Clk_period;
		Addr <=  "0100100010010";
		Trees_din <= x"dcff6508";
		wait for Clk_period;
		Addr <=  "0100100010011";
		Trees_din <= x"79ff1d04";
		wait for Clk_period;
		Addr <=  "0100100010100";
		Trees_din <= x"00542495";
		wait for Clk_period;
		Addr <=  "0100100010101";
		Trees_din <= x"ff932495";
		wait for Clk_period;
		Addr <=  "0100100010110";
		Trees_din <= x"ed004704";
		wait for Clk_period;
		Addr <=  "0100100010111";
		Trees_din <= x"ff6d2495";
		wait for Clk_period;
		Addr <=  "0100100011000";
		Trees_din <= x"fffd2495";
		wait for Clk_period;
		Addr <=  "0100100011001";
		Trees_din <= x"004a2495";
		wait for Clk_period;
		Addr <=  "0100100011010";
		Trees_din <= x"3bff7c10";
		wait for Clk_period;
		Addr <=  "0100100011011";
		Trees_din <= x"63ffa508";
		wait for Clk_period;
		Addr <=  "0100100011100";
		Trees_din <= x"5dffd104";
		wait for Clk_period;
		Addr <=  "0100100011101";
		Trees_din <= x"007a2495";
		wait for Clk_period;
		Addr <=  "0100100011110";
		Trees_din <= x"ffe02495";
		wait for Clk_period;
		Addr <=  "0100100011111";
		Trees_din <= x"30000804";
		wait for Clk_period;
		Addr <=  "0100100100000";
		Trees_din <= x"ff9f2495";
		wait for Clk_period;
		Addr <=  "0100100100001";
		Trees_din <= x"000d2495";
		wait for Clk_period;
		Addr <=  "0100100100010";
		Trees_din <= x"7cff9204";
		wait for Clk_period;
		Addr <=  "0100100100011";
		Trees_din <= x"ff932495";
		wait for Clk_period;
		Addr <=  "0100100100100";
		Trees_din <= x"ffea2495";
		wait for Clk_period;
		Addr <=  "0100100100101";
		Trees_din <= x"b8ff4564";
		wait for Clk_period;
		Addr <=  "0100100100110";
		Trees_din <= x"d9ff8f28";
		wait for Clk_period;
		Addr <=  "0100100100111";
		Trees_din <= x"bcff331c";
		wait for Clk_period;
		Addr <=  "0100100101000";
		Trees_din <= x"f8009d10";
		wait for Clk_period;
		Addr <=  "0100100101001";
		Trees_din <= x"71ff9f08";
		wait for Clk_period;
		Addr <=  "0100100101010";
		Trees_din <= x"1f012c04";
		wait for Clk_period;
		Addr <=  "0100100101011";
		Trees_din <= x"ffa52631";
		wait for Clk_period;
		Addr <=  "0100100101100";
		Trees_din <= x"00432631";
		wait for Clk_period;
		Addr <=  "0100100101101";
		Trees_din <= x"f1ffca04";
		wait for Clk_period;
		Addr <=  "0100100101110";
		Trees_din <= x"00732631";
		wait for Clk_period;
		Addr <=  "0100100101111";
		Trees_din <= x"ffd02631";
		wait for Clk_period;
		Addr <=  "0100100110000";
		Trees_din <= x"7fff5b08";
		wait for Clk_period;
		Addr <=  "0100100110001";
		Trees_din <= x"3bffa004";
		wait for Clk_period;
		Addr <=  "0100100110010";
		Trees_din <= x"ffa72631";
		wait for Clk_period;
		Addr <=  "0100100110011";
		Trees_din <= x"00322631";
		wait for Clk_period;
		Addr <=  "0100100110100";
		Trees_din <= x"00b32631";
		wait for Clk_period;
		Addr <=  "0100100110101";
		Trees_din <= x"ebff8708";
		wait for Clk_period;
		Addr <=  "0100100110110";
		Trees_din <= x"ddfe9c04";
		wait for Clk_period;
		Addr <=  "0100100110111";
		Trees_din <= x"001e2631";
		wait for Clk_period;
		Addr <=  "0100100111000";
		Trees_din <= x"ff6f2631";
		wait for Clk_period;
		Addr <=  "0100100111001";
		Trees_din <= x"00492631";
		wait for Clk_period;
		Addr <=  "0100100111010";
		Trees_din <= x"81ff751c";
		wait for Clk_period;
		Addr <=  "0100100111011";
		Trees_din <= x"34003c10";
		wait for Clk_period;
		Addr <=  "0100100111100";
		Trees_din <= x"e5fea308";
		wait for Clk_period;
		Addr <=  "0100100111101";
		Trees_din <= x"5ffefa04";
		wait for Clk_period;
		Addr <=  "0100100111110";
		Trees_din <= x"ff9c2631";
		wait for Clk_period;
		Addr <=  "0100100111111";
		Trees_din <= x"00342631";
		wait for Clk_period;
		Addr <=  "0100101000000";
		Trees_din <= x"ebff4504";
		wait for Clk_period;
		Addr <=  "0100101000001";
		Trees_din <= x"ff812631";
		wait for Clk_period;
		Addr <=  "0100101000010";
		Trees_din <= x"00002631";
		wait for Clk_period;
		Addr <=  "0100101000011";
		Trees_din <= x"ceffa408";
		wait for Clk_period;
		Addr <=  "0100101000100";
		Trees_din <= x"7cffc904";
		wait for Clk_period;
		Addr <=  "0100101000101";
		Trees_din <= x"00a32631";
		wait for Clk_period;
		Addr <=  "0100101000110";
		Trees_din <= x"00102631";
		wait for Clk_period;
		Addr <=  "0100101000111";
		Trees_din <= x"ffba2631";
		wait for Clk_period;
		Addr <=  "0100101001000";
		Trees_din <= x"efff1310";
		wait for Clk_period;
		Addr <=  "0100101001001";
		Trees_din <= x"d1ff3c08";
		wait for Clk_period;
		Addr <=  "0100101001010";
		Trees_din <= x"cb000804";
		wait for Clk_period;
		Addr <=  "0100101001011";
		Trees_din <= x"00af2631";
		wait for Clk_period;
		Addr <=  "0100101001100";
		Trees_din <= x"000b2631";
		wait for Clk_period;
		Addr <=  "0100101001101";
		Trees_din <= x"3f004e04";
		wait for Clk_period;
		Addr <=  "0100101001110";
		Trees_din <= x"ffab2631";
		wait for Clk_period;
		Addr <=  "0100101001111";
		Trees_din <= x"00732631";
		wait for Clk_period;
		Addr <=  "0100101010000";
		Trees_din <= x"a8ff8408";
		wait for Clk_period;
		Addr <=  "0100101010001";
		Trees_din <= x"bdffd204";
		wait for Clk_period;
		Addr <=  "0100101010010";
		Trees_din <= x"00572631";
		wait for Clk_period;
		Addr <=  "0100101010011";
		Trees_din <= x"fffc2631";
		wait for Clk_period;
		Addr <=  "0100101010100";
		Trees_din <= x"9dffa604";
		wait for Clk_period;
		Addr <=  "0100101010101";
		Trees_din <= x"ff942631";
		wait for Clk_period;
		Addr <=  "0100101010110";
		Trees_din <= x"00222631";
		wait for Clk_period;
		Addr <=  "0100101010111";
		Trees_din <= x"26001d30";
		wait for Clk_period;
		Addr <=  "0100101011000";
		Trees_din <= x"a4ff7518";
		wait for Clk_period;
		Addr <=  "0100101011001";
		Trees_din <= x"e1ff9308";
		wait for Clk_period;
		Addr <=  "0100101011010";
		Trees_din <= x"f1ffe104";
		wait for Clk_period;
		Addr <=  "0100101011011";
		Trees_din <= x"ff7e2631";
		wait for Clk_period;
		Addr <=  "0100101011100";
		Trees_din <= x"ffdd2631";
		wait for Clk_period;
		Addr <=  "0100101011101";
		Trees_din <= x"6e001008";
		wait for Clk_period;
		Addr <=  "0100101011110";
		Trees_din <= x"30005f04";
		wait for Clk_period;
		Addr <=  "0100101011111";
		Trees_din <= x"ff842631";
		wait for Clk_period;
		Addr <=  "0100101100000";
		Trees_din <= x"00422631";
		wait for Clk_period;
		Addr <=  "0100101100001";
		Trees_din <= x"a9ff6b04";
		wait for Clk_period;
		Addr <=  "0100101100010";
		Trees_din <= x"00792631";
		wait for Clk_period;
		Addr <=  "0100101100011";
		Trees_din <= x"ffdd2631";
		wait for Clk_period;
		Addr <=  "0100101100100";
		Trees_din <= x"65fef90c";
		wait for Clk_period;
		Addr <=  "0100101100101";
		Trees_din <= x"c8005008";
		wait for Clk_period;
		Addr <=  "0100101100110";
		Trees_din <= x"34ffea04";
		wait for Clk_period;
		Addr <=  "0100101100111";
		Trees_din <= x"00052631";
		wait for Clk_period;
		Addr <=  "0100101101000";
		Trees_din <= x"ff952631";
		wait for Clk_period;
		Addr <=  "0100101101001";
		Trees_din <= x"00792631";
		wait for Clk_period;
		Addr <=  "0100101101010";
		Trees_din <= x"dc008f08";
		wait for Clk_period;
		Addr <=  "0100101101011";
		Trees_din <= x"b8ff5404";
		wait for Clk_period;
		Addr <=  "0100101101100";
		Trees_din <= x"fffe2631";
		wait for Clk_period;
		Addr <=  "0100101101101";
		Trees_din <= x"ff702631";
		wait for Clk_period;
		Addr <=  "0100101101110";
		Trees_din <= x"001f2631";
		wait for Clk_period;
		Addr <=  "0100101101111";
		Trees_din <= x"a2ffa61c";
		wait for Clk_period;
		Addr <=  "0100101110000";
		Trees_din <= x"24fff110";
		wait for Clk_period;
		Addr <=  "0100101110001";
		Trees_din <= x"64ff4108";
		wait for Clk_period;
		Addr <=  "0100101110010";
		Trees_din <= x"6d005704";
		wait for Clk_period;
		Addr <=  "0100101110011";
		Trees_din <= x"003f2631";
		wait for Clk_period;
		Addr <=  "0100101110100";
		Trees_din <= x"ffba2631";
		wait for Clk_period;
		Addr <=  "0100101110101";
		Trees_din <= x"74000a04";
		wait for Clk_period;
		Addr <=  "0100101110110";
		Trees_din <= x"ff8f2631";
		wait for Clk_period;
		Addr <=  "0100101110111";
		Trees_din <= x"00082631";
		wait for Clk_period;
		Addr <=  "0100101111000";
		Trees_din <= x"5eff4104";
		wait for Clk_period;
		Addr <=  "0100101111001";
		Trees_din <= x"ffa02631";
		wait for Clk_period;
		Addr <=  "0100101111010";
		Trees_din <= x"6effe204";
		wait for Clk_period;
		Addr <=  "0100101111011";
		Trees_din <= x"ffc32631";
		wait for Clk_period;
		Addr <=  "0100101111100";
		Trees_din <= x"00812631";
		wait for Clk_period;
		Addr <=  "0100101111101";
		Trees_din <= x"f6fed610";
		wait for Clk_period;
		Addr <=  "0100101111110";
		Trees_din <= x"20007708";
		wait for Clk_period;
		Addr <=  "0100101111111";
		Trees_din <= x"77ff7404";
		wait for Clk_period;
		Addr <=  "0100110000000";
		Trees_din <= x"ff922631";
		wait for Clk_period;
		Addr <=  "0100110000001";
		Trees_din <= x"00082631";
		wait for Clk_period;
		Addr <=  "0100110000010";
		Trees_din <= x"22006804";
		wait for Clk_period;
		Addr <=  "0100110000011";
		Trees_din <= x"00182631";
		wait for Clk_period;
		Addr <=  "0100110000100";
		Trees_din <= x"00812631";
		wait for Clk_period;
		Addr <=  "0100110000101";
		Trees_din <= x"1fffa308";
		wait for Clk_period;
		Addr <=  "0100110000110";
		Trees_din <= x"f7ff5104";
		wait for Clk_period;
		Addr <=  "0100110000111";
		Trees_din <= x"005d2631";
		wait for Clk_period;
		Addr <=  "0100110001000";
		Trees_din <= x"fff32631";
		wait for Clk_period;
		Addr <=  "0100110001001";
		Trees_din <= x"2effbe04";
		wait for Clk_period;
		Addr <=  "0100110001010";
		Trees_din <= x"ffb22631";
		wait for Clk_period;
		Addr <=  "0100110001011";
		Trees_din <= x"000d2631";
		wait for Clk_period;
		Addr <=  "0100110001100";
		Trees_din <= x"01fe7b4c";
		wait for Clk_period;
		Addr <=  "0100110001101";
		Trees_din <= x"2cff1a10";
		wait for Clk_period;
		Addr <=  "0100110001110";
		Trees_din <= x"3aff1504";
		wait for Clk_period;
		Addr <=  "0100110001111";
		Trees_din <= x"ff7c27b5";
		wait for Clk_period;
		Addr <=  "0100110010000";
		Trees_din <= x"9bff1b08";
		wait for Clk_period;
		Addr <=  "0100110010001";
		Trees_din <= x"d3ff0304";
		wait for Clk_period;
		Addr <=  "0100110010010";
		Trees_din <= x"ffcf27b5";
		wait for Clk_period;
		Addr <=  "0100110010011";
		Trees_din <= x"007a27b5";
		wait for Clk_period;
		Addr <=  "0100110010100";
		Trees_din <= x"ffb127b5";
		wait for Clk_period;
		Addr <=  "0100110010101";
		Trees_din <= x"be004020";
		wait for Clk_period;
		Addr <=  "0100110010110";
		Trees_din <= x"edffc210";
		wait for Clk_period;
		Addr <=  "0100110010111";
		Trees_din <= x"34000708";
		wait for Clk_period;
		Addr <=  "0100110011000";
		Trees_din <= x"87ff7004";
		wait for Clk_period;
		Addr <=  "0100110011001";
		Trees_din <= x"ffdf27b5";
		wait for Clk_period;
		Addr <=  "0100110011010";
		Trees_din <= x"005027b5";
		wait for Clk_period;
		Addr <=  "0100110011011";
		Trees_din <= x"cafd8404";
		wait for Clk_period;
		Addr <=  "0100110011100";
		Trees_din <= x"003e27b5";
		wait for Clk_period;
		Addr <=  "0100110011101";
		Trees_din <= x"ffab27b5";
		wait for Clk_period;
		Addr <=  "0100110011110";
		Trees_din <= x"9a001508";
		wait for Clk_period;
		Addr <=  "0100110011111";
		Trees_din <= x"58ff7504";
		wait for Clk_period;
		Addr <=  "0100110100000";
		Trees_din <= x"004727b5";
		wait for Clk_period;
		Addr <=  "0100110100001";
		Trees_din <= x"ffc227b5";
		wait for Clk_period;
		Addr <=  "0100110100010";
		Trees_din <= x"90ff8f04";
		wait for Clk_period;
		Addr <=  "0100110100011";
		Trees_din <= x"ff8727b5";
		wait for Clk_period;
		Addr <=  "0100110100100";
		Trees_din <= x"003127b5";
		wait for Clk_period;
		Addr <=  "0100110100101";
		Trees_din <= x"53ff5a0c";
		wait for Clk_period;
		Addr <=  "0100110100110";
		Trees_din <= x"35fe7b04";
		wait for Clk_period;
		Addr <=  "0100110100111";
		Trees_din <= x"ffea27b5";
		wait for Clk_period;
		Addr <=  "0100110101000";
		Trees_din <= x"6bfeea04";
		wait for Clk_period;
		Addr <=  "0100110101001";
		Trees_din <= x"004427b5";
		wait for Clk_period;
		Addr <=  "0100110101010";
		Trees_din <= x"00b827b5";
		wait for Clk_period;
		Addr <=  "0100110101011";
		Trees_din <= x"bbfef708";
		wait for Clk_period;
		Addr <=  "0100110101100";
		Trees_din <= x"5fff6a04";
		wait for Clk_period;
		Addr <=  "0100110101101";
		Trees_din <= x"ff8c27b5";
		wait for Clk_period;
		Addr <=  "0100110101110";
		Trees_din <= x"003027b5";
		wait for Clk_period;
		Addr <=  "0100110101111";
		Trees_din <= x"72000a04";
		wait for Clk_period;
		Addr <=  "0100110110000";
		Trees_din <= x"007927b5";
		wait for Clk_period;
		Addr <=  "0100110110001";
		Trees_din <= x"001027b5";
		wait for Clk_period;
		Addr <=  "0100110110010";
		Trees_din <= x"fbff8b3c";
		wait for Clk_period;
		Addr <=  "0100110110011";
		Trees_din <= x"f1ffad1c";
		wait for Clk_period;
		Addr <=  "0100110110100";
		Trees_din <= x"8cfffb10";
		wait for Clk_period;
		Addr <=  "0100110110101";
		Trees_din <= x"3eff5f08";
		wait for Clk_period;
		Addr <=  "0100110110110";
		Trees_din <= x"72000604";
		wait for Clk_period;
		Addr <=  "0100110110111";
		Trees_din <= x"ffc527b5";
		wait for Clk_period;
		Addr <=  "0100110111000";
		Trees_din <= x"006527b5";
		wait for Clk_period;
		Addr <=  "0100110111001";
		Trees_din <= x"62ff0e04";
		wait for Clk_period;
		Addr <=  "0100110111010";
		Trees_din <= x"002b27b5";
		wait for Clk_period;
		Addr <=  "0100110111011";
		Trees_din <= x"ffa927b5";
		wait for Clk_period;
		Addr <=  "0100110111100";
		Trees_din <= x"2fff1904";
		wait for Clk_period;
		Addr <=  "0100110111101";
		Trees_din <= x"ffa227b5";
		wait for Clk_period;
		Addr <=  "0100110111110";
		Trees_din <= x"85ff4c04";
		wait for Clk_period;
		Addr <=  "0100110111111";
		Trees_din <= x"000027b5";
		wait for Clk_period;
		Addr <=  "0100111000000";
		Trees_din <= x"00a327b5";
		wait for Clk_period;
		Addr <=  "0100111000001";
		Trees_din <= x"34002310";
		wait for Clk_period;
		Addr <=  "0100111000010";
		Trees_din <= x"b3ff6b08";
		wait for Clk_period;
		Addr <=  "0100111000011";
		Trees_din <= x"8dff8004";
		wait for Clk_period;
		Addr <=  "0100111000100";
		Trees_din <= x"ff9f27b5";
		wait for Clk_period;
		Addr <=  "0100111000101";
		Trees_din <= x"003127b5";
		wait for Clk_period;
		Addr <=  "0100111000110";
		Trees_din <= x"b6ff2c04";
		wait for Clk_period;
		Addr <=  "0100111000111";
		Trees_din <= x"ffa927b5";
		wait for Clk_period;
		Addr <=  "0100111001000";
		Trees_din <= x"005f27b5";
		wait for Clk_period;
		Addr <=  "0100111001001";
		Trees_din <= x"87ff7008";
		wait for Clk_period;
		Addr <=  "0100111001010";
		Trees_din <= x"e8ffe204";
		wait for Clk_period;
		Addr <=  "0100111001011";
		Trees_din <= x"ff9127b5";
		wait for Clk_period;
		Addr <=  "0100111001100";
		Trees_din <= x"003727b5";
		wait for Clk_period;
		Addr <=  "0100111001101";
		Trees_din <= x"56ff8904";
		wait for Clk_period;
		Addr <=  "0100111001110";
		Trees_din <= x"008227b5";
		wait for Clk_period;
		Addr <=  "0100111001111";
		Trees_din <= x"ffcd27b5";
		wait for Clk_period;
		Addr <=  "0100111010000";
		Trees_din <= x"45fec81c";
		wait for Clk_period;
		Addr <=  "0100111010001";
		Trees_din <= x"90001b10";
		wait for Clk_period;
		Addr <=  "0100111010010";
		Trees_din <= x"d9001208";
		wait for Clk_period;
		Addr <=  "0100111010011";
		Trees_din <= x"ee009004";
		wait for Clk_period;
		Addr <=  "0100111010100";
		Trees_din <= x"ff8327b5";
		wait for Clk_period;
		Addr <=  "0100111010101";
		Trees_din <= x"001027b5";
		wait for Clk_period;
		Addr <=  "0100111010110";
		Trees_din <= x"1effd004";
		wait for Clk_period;
		Addr <=  "0100111010111";
		Trees_din <= x"ff9c27b5";
		wait for Clk_period;
		Addr <=  "0100111011000";
		Trees_din <= x"005a27b5";
		wait for Clk_period;
		Addr <=  "0100111011001";
		Trees_din <= x"cafe7708";
		wait for Clk_period;
		Addr <=  "0100111011010";
		Trees_din <= x"36ff4a04";
		wait for Clk_period;
		Addr <=  "0100111011011";
		Trees_din <= x"009527b5";
		wait for Clk_period;
		Addr <=  "0100111011100";
		Trees_din <= x"ffe827b5";
		wait for Clk_period;
		Addr <=  "0100111011101";
		Trees_din <= x"ffab27b5";
		wait for Clk_period;
		Addr <=  "0100111011110";
		Trees_din <= x"86ff1d10";
		wait for Clk_period;
		Addr <=  "0100111011111";
		Trees_din <= x"28ff0508";
		wait for Clk_period;
		Addr <=  "0100111100000";
		Trees_din <= x"0efee604";
		wait for Clk_period;
		Addr <=  "0100111100001";
		Trees_din <= x"004f27b5";
		wait for Clk_period;
		Addr <=  "0100111100010";
		Trees_din <= x"ff9d27b5";
		wait for Clk_period;
		Addr <=  "0100111100011";
		Trees_din <= x"17006104";
		wait for Clk_period;
		Addr <=  "0100111100100";
		Trees_din <= x"ff8327b5";
		wait for Clk_period;
		Addr <=  "0100111100101";
		Trees_din <= x"001127b5";
		wait for Clk_period;
		Addr <=  "0100111100110";
		Trees_din <= x"55002108";
		wait for Clk_period;
		Addr <=  "0100111100111";
		Trees_din <= x"6d002b04";
		wait for Clk_period;
		Addr <=  "0100111101000";
		Trees_din <= x"ff9927b5";
		wait for Clk_period;
		Addr <=  "0100111101001";
		Trees_din <= x"001a27b5";
		wait for Clk_period;
		Addr <=  "0100111101010";
		Trees_din <= x"41fef104";
		wait for Clk_period;
		Addr <=  "0100111101011";
		Trees_din <= x"ffe827b5";
		wait for Clk_period;
		Addr <=  "0100111101100";
		Trees_din <= x"005727b5";
		wait for Clk_period;
		Addr <=  "0100111101101";
		Trees_din <= x"cbff392c";
		wait for Clk_period;
		Addr <=  "0100111101110";
		Trees_din <= x"4effc620";
		wait for Clk_period;
		Addr <=  "0100111101111";
		Trees_din <= x"a6ffa810";
		wait for Clk_period;
		Addr <=  "0100111110000";
		Trees_din <= x"0701190c";
		wait for Clk_period;
		Addr <=  "0100111110001";
		Trees_din <= x"79fed404";
		wait for Clk_period;
		Addr <=  "0100111110010";
		Trees_din <= x"002328e1";
		wait for Clk_period;
		Addr <=  "0100111110011";
		Trees_din <= x"ccff0e04";
		wait for Clk_period;
		Addr <=  "0100111110100";
		Trees_din <= x"ffec28e1";
		wait for Clk_period;
		Addr <=  "0100111110101";
		Trees_din <= x"ff6a28e1";
		wait for Clk_period;
		Addr <=  "0100111110110";
		Trees_din <= x"002428e1";
		wait for Clk_period;
		Addr <=  "0100111110111";
		Trees_din <= x"24ffca08";
		wait for Clk_period;
		Addr <=  "0100111111000";
		Trees_din <= x"70fe9604";
		wait for Clk_period;
		Addr <=  "0100111111001";
		Trees_din <= x"002128e1";
		wait for Clk_period;
		Addr <=  "0100111111010";
		Trees_din <= x"ff8e28e1";
		wait for Clk_period;
		Addr <=  "0100111111011";
		Trees_din <= x"f6ff3704";
		wait for Clk_period;
		Addr <=  "0100111111100";
		Trees_din <= x"000b28e1";
		wait for Clk_period;
		Addr <=  "0100111111101";
		Trees_din <= x"009928e1";
		wait for Clk_period;
		Addr <=  "0100111111110";
		Trees_din <= x"3eff8108";
		wait for Clk_period;
		Addr <=  "0100111111111";
		Trees_din <= x"3f001804";
		wait for Clk_period;
		Addr <=  "0101000000000";
		Trees_din <= x"fff028e1";
		wait for Clk_period;
		Addr <=  "0101000000001";
		Trees_din <= x"008c28e1";
		wait for Clk_period;
		Addr <=  "0101000000010";
		Trees_din <= x"ffbe28e1";
		wait for Clk_period;
		Addr <=  "0101000000011";
		Trees_din <= x"c7fea030";
		wait for Clk_period;
		Addr <=  "0101000000100";
		Trees_din <= x"87ff8818";
		wait for Clk_period;
		Addr <=  "0101000000101";
		Trees_din <= x"5d000710";
		wait for Clk_period;
		Addr <=  "0101000000110";
		Trees_din <= x"54009d08";
		wait for Clk_period;
		Addr <=  "0101000000111";
		Trees_din <= x"ce002504";
		wait for Clk_period;
		Addr <=  "0101000001000";
		Trees_din <= x"002f28e1";
		wait for Clk_period;
		Addr <=  "0101000001001";
		Trees_din <= x"ffb928e1";
		wait for Clk_period;
		Addr <=  "0101000001010";
		Trees_din <= x"ceff2804";
		wait for Clk_period;
		Addr <=  "0101000001011";
		Trees_din <= x"006a28e1";
		wait for Clk_period;
		Addr <=  "0101000001100";
		Trees_din <= x"ff9c28e1";
		wait for Clk_period;
		Addr <=  "0101000001101";
		Trees_din <= x"fcffab04";
		wait for Clk_period;
		Addr <=  "0101000001110";
		Trees_din <= x"ff8228e1";
		wait for Clk_period;
		Addr <=  "0101000001111";
		Trees_din <= x"000c28e1";
		wait for Clk_period;
		Addr <=  "0101000010000";
		Trees_din <= x"42fed208";
		wait for Clk_period;
		Addr <=  "0101000010001";
		Trees_din <= x"7affed04";
		wait for Clk_period;
		Addr <=  "0101000010010";
		Trees_din <= x"ffd328e1";
		wait for Clk_period;
		Addr <=  "0101000010011";
		Trees_din <= x"006828e1";
		wait for Clk_period;
		Addr <=  "0101000010100";
		Trees_din <= x"05002008";
		wait for Clk_period;
		Addr <=  "0101000010101";
		Trees_din <= x"04009404";
		wait for Clk_period;
		Addr <=  "0101000010110";
		Trees_din <= x"ffb028e1";
		wait for Clk_period;
		Addr <=  "0101000010111";
		Trees_din <= x"006128e1";
		wait for Clk_period;
		Addr <=  "0101000011000";
		Trees_din <= x"56fe8c04";
		wait for Clk_period;
		Addr <=  "0101000011001";
		Trees_din <= x"000528e1";
		wait for Clk_period;
		Addr <=  "0101000011010";
		Trees_din <= x"ff7128e1";
		wait for Clk_period;
		Addr <=  "0101000011011";
		Trees_din <= x"b8ff4520";
		wait for Clk_period;
		Addr <=  "0101000011100";
		Trees_din <= x"d9ff8410";
		wait for Clk_period;
		Addr <=  "0101000011101";
		Trees_din <= x"40003008";
		wait for Clk_period;
		Addr <=  "0101000011110";
		Trees_din <= x"ddff9004";
		wait for Clk_period;
		Addr <=  "0101000011111";
		Trees_din <= x"ff8428e1";
		wait for Clk_period;
		Addr <=  "0101000100000";
		Trees_din <= x"001228e1";
		wait for Clk_period;
		Addr <=  "0101000100001";
		Trees_din <= x"33feff04";
		wait for Clk_period;
		Addr <=  "0101000100010";
		Trees_din <= x"ffb528e1";
		wait for Clk_period;
		Addr <=  "0101000100011";
		Trees_din <= x"005f28e1";
		wait for Clk_period;
		Addr <=  "0101000100100";
		Trees_din <= x"d8007a08";
		wait for Clk_period;
		Addr <=  "0101000100101";
		Trees_din <= x"ebff2504";
		wait for Clk_period;
		Addr <=  "0101000100110";
		Trees_din <= x"005528e1";
		wait for Clk_period;
		Addr <=  "0101000100111";
		Trees_din <= x"fffa28e1";
		wait for Clk_period;
		Addr <=  "0101000101000";
		Trees_din <= x"72007604";
		wait for Clk_period;
		Addr <=  "0101000101001";
		Trees_din <= x"ffb528e1";
		wait for Clk_period;
		Addr <=  "0101000101010";
		Trees_din <= x"004f28e1";
		wait for Clk_period;
		Addr <=  "0101000101011";
		Trees_din <= x"cfff8e0c";
		wait for Clk_period;
		Addr <=  "0101000101100";
		Trees_din <= x"b3ff0404";
		wait for Clk_period;
		Addr <=  "0101000101101";
		Trees_din <= x"ffa828e1";
		wait for Clk_period;
		Addr <=  "0101000101110";
		Trees_din <= x"76ff7104";
		wait for Clk_period;
		Addr <=  "0101000101111";
		Trees_din <= x"ffc728e1";
		wait for Clk_period;
		Addr <=  "0101000110000";
		Trees_din <= x"008028e1";
		wait for Clk_period;
		Addr <=  "0101000110001";
		Trees_din <= x"5a007a08";
		wait for Clk_period;
		Addr <=  "0101000110010";
		Trees_din <= x"daffbf04";
		wait for Clk_period;
		Addr <=  "0101000110011";
		Trees_din <= x"002f28e1";
		wait for Clk_period;
		Addr <=  "0101000110100";
		Trees_din <= x"fff028e1";
		wait for Clk_period;
		Addr <=  "0101000110101";
		Trees_din <= x"50ffb104";
		wait for Clk_period;
		Addr <=  "0101000110110";
		Trees_din <= x"ffbb28e1";
		wait for Clk_period;
		Addr <=  "0101000110111";
		Trees_din <= x"002428e1";
		wait for Clk_period;
		Addr <=  "0101000111000";
		Trees_din <= x"6f003e54";
		wait for Clk_period;
		Addr <=  "0101000111001";
		Trees_din <= x"feff992c";
		wait for Clk_period;
		Addr <=  "0101000111010";
		Trees_din <= x"a5ff6720";
		wait for Clk_period;
		Addr <=  "0101000111011";
		Trees_din <= x"be001910";
		wait for Clk_period;
		Addr <=  "0101000111100";
		Trees_din <= x"a4ff5108";
		wait for Clk_period;
		Addr <=  "0101000111101";
		Trees_din <= x"17ffe204";
		wait for Clk_period;
		Addr <=  "0101000111110";
		Trees_din <= x"ffcc299d";
		wait for Clk_period;
		Addr <=  "0101000111111";
		Trees_din <= x"0042299d";
		wait for Clk_period;
		Addr <=  "0101001000000";
		Trees_din <= x"0efe1104";
		wait for Clk_period;
		Addr <=  "0101001000001";
		Trees_din <= x"0027299d";
		wait for Clk_period;
		Addr <=  "0101001000010";
		Trees_din <= x"ffb5299d";
		wait for Clk_period;
		Addr <=  "0101001000011";
		Trees_din <= x"fdff9808";
		wait for Clk_period;
		Addr <=  "0101001000100";
		Trees_din <= x"49ffe904";
		wait for Clk_period;
		Addr <=  "0101001000101";
		Trees_din <= x"fff9299d";
		wait for Clk_period;
		Addr <=  "0101001000110";
		Trees_din <= x"0042299d";
		wait for Clk_period;
		Addr <=  "0101001000111";
		Trees_din <= x"a5fecf04";
		wait for Clk_period;
		Addr <=  "0101001001000";
		Trees_din <= x"0037299d";
		wait for Clk_period;
		Addr <=  "0101001001001";
		Trees_din <= x"ff93299d";
		wait for Clk_period;
		Addr <=  "0101001001010";
		Trees_din <= x"cafd9004";
		wait for Clk_period;
		Addr <=  "0101001001011";
		Trees_din <= x"0046299d";
		wait for Clk_period;
		Addr <=  "0101001001100";
		Trees_din <= x"aefe3b04";
		wait for Clk_period;
		Addr <=  "0101001001101";
		Trees_din <= x"0016299d";
		wait for Clk_period;
		Addr <=  "0101001001110";
		Trees_din <= x"ff73299d";
		wait for Clk_period;
		Addr <=  "0101001001111";
		Trees_din <= x"44ff5608";
		wait for Clk_period;
		Addr <=  "0101001010000";
		Trees_din <= x"64fecd04";
		wait for Clk_period;
		Addr <=  "0101001010001";
		Trees_din <= x"000f299d";
		wait for Clk_period;
		Addr <=  "0101001010010";
		Trees_din <= x"ff7c299d";
		wait for Clk_period;
		Addr <=  "0101001010011";
		Trees_din <= x"c3001610";
		wait for Clk_period;
		Addr <=  "0101001010100";
		Trees_din <= x"01fef708";
		wait for Clk_period;
		Addr <=  "0101001010101";
		Trees_din <= x"bffe8a04";
		wait for Clk_period;
		Addr <=  "0101001010110";
		Trees_din <= x"ffca299d";
		wait for Clk_period;
		Addr <=  "0101001010111";
		Trees_din <= x"0037299d";
		wait for Clk_period;
		Addr <=  "0101001011000";
		Trees_din <= x"dafff504";
		wait for Clk_period;
		Addr <=  "0101001011001";
		Trees_din <= x"ffad299d";
		wait for Clk_period;
		Addr <=  "0101001011010";
		Trees_din <= x"001f299d";
		wait for Clk_period;
		Addr <=  "0101001011011";
		Trees_din <= x"ddfeef08";
		wait for Clk_period;
		Addr <=  "0101001011100";
		Trees_din <= x"cfffd204";
		wait for Clk_period;
		Addr <=  "0101001011101";
		Trees_din <= x"0091299d";
		wait for Clk_period;
		Addr <=  "0101001011110";
		Trees_din <= x"fffb299d";
		wait for Clk_period;
		Addr <=  "0101001011111";
		Trees_din <= x"45fecf04";
		wait for Clk_period;
		Addr <=  "0101001100000";
		Trees_din <= x"ff95299d";
		wait for Clk_period;
		Addr <=  "0101001100001";
		Trees_din <= x"fff9299d";
		wait for Clk_period;
		Addr <=  "0101001100010";
		Trees_din <= x"3eff1a04";
		wait for Clk_period;
		Addr <=  "0101001100011";
		Trees_din <= x"0026299d";
		wait for Clk_period;
		Addr <=  "0101001100100";
		Trees_din <= x"0b007404";
		wait for Clk_period;
		Addr <=  "0101001100101";
		Trees_din <= x"ff7e299d";
		wait for Clk_period;
		Addr <=  "0101001100110";
		Trees_din <= x"ffee299d";
		wait for Clk_period;
		Addr <=  "0101001100111";
		Trees_din <= x"69feb928";
		wait for Clk_period;
		Addr <=  "0101001101000";
		Trees_din <= x"55ffcb10";
		wait for Clk_period;
		Addr <=  "0101001101001";
		Trees_din <= x"75003104";
		wait for Clk_period;
		Addr <=  "0101001101010";
		Trees_din <= x"ff972a91";
		wait for Clk_period;
		Addr <=  "0101001101011";
		Trees_din <= x"48ff4c04";
		wait for Clk_period;
		Addr <=  "0101001101100";
		Trees_din <= x"ffa82a91";
		wait for Clk_period;
		Addr <=  "0101001101101";
		Trees_din <= x"b7ff7e04";
		wait for Clk_period;
		Addr <=  "0101001101110";
		Trees_din <= x"00662a91";
		wait for Clk_period;
		Addr <=  "0101001101111";
		Trees_din <= x"fff02a91";
		wait for Clk_period;
		Addr <=  "0101001110000";
		Trees_din <= x"71ffe414";
		wait for Clk_period;
		Addr <=  "0101001110001";
		Trees_din <= x"bbffde10";
		wait for Clk_period;
		Addr <=  "0101001110010";
		Trees_din <= x"6bfe9b08";
		wait for Clk_period;
		Addr <=  "0101001110011";
		Trees_din <= x"64fef004";
		wait for Clk_period;
		Addr <=  "0101001110100";
		Trees_din <= x"004d2a91";
		wait for Clk_period;
		Addr <=  "0101001110101";
		Trees_din <= x"ffd62a91";
		wait for Clk_period;
		Addr <=  "0101001110110";
		Trees_din <= x"22ff7b04";
		wait for Clk_period;
		Addr <=  "0101001110111";
		Trees_din <= x"ffed2a91";
		wait for Clk_period;
		Addr <=  "0101001111000";
		Trees_din <= x"00772a91";
		wait for Clk_period;
		Addr <=  "0101001111001";
		Trees_din <= x"ffbe2a91";
		wait for Clk_period;
		Addr <=  "0101001111010";
		Trees_din <= x"ffaa2a91";
		wait for Clk_period;
		Addr <=  "0101001111011";
		Trees_din <= x"5eff2b14";
		wait for Clk_period;
		Addr <=  "0101001111100";
		Trees_din <= x"b5ff620c";
		wait for Clk_period;
		Addr <=  "0101001111101";
		Trees_din <= x"4700b108";
		wait for Clk_period;
		Addr <=  "0101001111110";
		Trees_din <= x"f9fe6d04";
		wait for Clk_period;
		Addr <=  "0101001111111";
		Trees_din <= x"ffd92a91";
		wait for Clk_period;
		Addr <=  "0101010000000";
		Trees_din <= x"ff732a91";
		wait for Clk_period;
		Addr <=  "0101010000001";
		Trees_din <= x"00292a91";
		wait for Clk_period;
		Addr <=  "0101010000010";
		Trees_din <= x"76ff9204";
		wait for Clk_period;
		Addr <=  "0101010000011";
		Trees_din <= x"00692a91";
		wait for Clk_period;
		Addr <=  "0101010000100";
		Trees_din <= x"ffe32a91";
		wait for Clk_period;
		Addr <=  "0101010000101";
		Trees_din <= x"76ffc920";
		wait for Clk_period;
		Addr <=  "0101010000110";
		Trees_din <= x"29ffc110";
		wait for Clk_period;
		Addr <=  "0101010000111";
		Trees_din <= x"ee009208";
		wait for Clk_period;
		Addr <=  "0101010001000";
		Trees_din <= x"70ff0c04";
		wait for Clk_period;
		Addr <=  "0101010001001";
		Trees_din <= x"ffde2a91";
		wait for Clk_period;
		Addr <=  "0101010001010";
		Trees_din <= x"00152a91";
		wait for Clk_period;
		Addr <=  "0101010001011";
		Trees_din <= x"eaff6504";
		wait for Clk_period;
		Addr <=  "0101010001100";
		Trees_din <= x"ffc82a91";
		wait for Clk_period;
		Addr <=  "0101010001101";
		Trees_din <= x"007b2a91";
		wait for Clk_period;
		Addr <=  "0101010001110";
		Trees_din <= x"d5002e08";
		wait for Clk_period;
		Addr <=  "0101010001111";
		Trees_din <= x"a3ffec04";
		wait for Clk_period;
		Addr <=  "0101010010000";
		Trees_din <= x"ff7a2a91";
		wait for Clk_period;
		Addr <=  "0101010010001";
		Trees_din <= x"00092a91";
		wait for Clk_period;
		Addr <=  "0101010010010";
		Trees_din <= x"16ff0604";
		wait for Clk_period;
		Addr <=  "0101010010011";
		Trees_din <= x"ffb92a91";
		wait for Clk_period;
		Addr <=  "0101010010100";
		Trees_din <= x"004b2a91";
		wait for Clk_period;
		Addr <=  "0101010010101";
		Trees_din <= x"07ffc810";
		wait for Clk_period;
		Addr <=  "0101010010110";
		Trees_din <= x"26ffee08";
		wait for Clk_period;
		Addr <=  "0101010010111";
		Trees_din <= x"f6fef704";
		wait for Clk_period;
		Addr <=  "0101010011000";
		Trees_din <= x"fffc2a91";
		wait for Clk_period;
		Addr <=  "0101010011001";
		Trees_din <= x"ffa62a91";
		wait for Clk_period;
		Addr <=  "0101010011010";
		Trees_din <= x"42ffde04";
		wait for Clk_period;
		Addr <=  "0101010011011";
		Trees_din <= x"00862a91";
		wait for Clk_period;
		Addr <=  "0101010011100";
		Trees_din <= x"ffc02a91";
		wait for Clk_period;
		Addr <=  "0101010011101";
		Trees_din <= x"ebfe6208";
		wait for Clk_period;
		Addr <=  "0101010011110";
		Trees_din <= x"9bfeee04";
		wait for Clk_period;
		Addr <=  "0101010011111";
		Trees_din <= x"fff02a91";
		wait for Clk_period;
		Addr <=  "0101010100000";
		Trees_din <= x"ff812a91";
		wait for Clk_period;
		Addr <=  "0101010100001";
		Trees_din <= x"ecff7d04";
		wait for Clk_period;
		Addr <=  "0101010100010";
		Trees_din <= x"ffb92a91";
		wait for Clk_period;
		Addr <=  "0101010100011";
		Trees_din <= x"00132a91";
		wait for Clk_period;
		Addr <=  "0101010100100";
		Trees_din <= x"e7ff7b4c";
		wait for Clk_period;
		Addr <=  "0101010100101";
		Trees_din <= x"20ff2e14";
		wait for Clk_period;
		Addr <=  "0101010100110";
		Trees_din <= x"fb001d0c";
		wait for Clk_period;
		Addr <=  "0101010100111";
		Trees_din <= x"9eff2408";
		wait for Clk_period;
		Addr <=  "0101010101000";
		Trees_din <= x"ab00ef04";
		wait for Clk_period;
		Addr <=  "0101010101001";
		Trees_din <= x"ffb52bd5";
		wait for Clk_period;
		Addr <=  "0101010101010";
		Trees_din <= x"003c2bd5";
		wait for Clk_period;
		Addr <=  "0101010101011";
		Trees_din <= x"ff792bd5";
		wait for Clk_period;
		Addr <=  "0101010101100";
		Trees_din <= x"2cff5c04";
		wait for Clk_period;
		Addr <=  "0101010101101";
		Trees_din <= x"007c2bd5";
		wait for Clk_period;
		Addr <=  "0101010101110";
		Trees_din <= x"ffc02bd5";
		wait for Clk_period;
		Addr <=  "0101010101111";
		Trees_din <= x"eaff3520";
		wait for Clk_period;
		Addr <=  "0101010110000";
		Trees_din <= x"30fff610";
		wait for Clk_period;
		Addr <=  "0101010110001";
		Trees_din <= x"e7ff0d08";
		wait for Clk_period;
		Addr <=  "0101010110010";
		Trees_din <= x"66ffd704";
		wait for Clk_period;
		Addr <=  "0101010110011";
		Trees_din <= x"004f2bd5";
		wait for Clk_period;
		Addr <=  "0101010110100";
		Trees_din <= x"ffb82bd5";
		wait for Clk_period;
		Addr <=  "0101010110101";
		Trees_din <= x"e3ff1404";
		wait for Clk_period;
		Addr <=  "0101010110110";
		Trees_din <= x"ff772bd5";
		wait for Clk_period;
		Addr <=  "0101010110111";
		Trees_din <= x"fff52bd5";
		wait for Clk_period;
		Addr <=  "0101010111000";
		Trees_din <= x"10ffe808";
		wait for Clk_period;
		Addr <=  "0101010111001";
		Trees_din <= x"7fff5304";
		wait for Clk_period;
		Addr <=  "0101010111010";
		Trees_din <= x"ffa22bd5";
		wait for Clk_period;
		Addr <=  "0101010111011";
		Trees_din <= x"00042bd5";
		wait for Clk_period;
		Addr <=  "0101010111100";
		Trees_din <= x"cf003004";
		wait for Clk_period;
		Addr <=  "0101010111101";
		Trees_din <= x"fffd2bd5";
		wait for Clk_period;
		Addr <=  "0101010111110";
		Trees_din <= x"007d2bd5";
		wait for Clk_period;
		Addr <=  "0101010111111";
		Trees_din <= x"5eff2e08";
		wait for Clk_period;
		Addr <=  "0101011000000";
		Trees_din <= x"a1fe9a04";
		wait for Clk_period;
		Addr <=  "0101011000001";
		Trees_din <= x"00122bd5";
		wait for Clk_period;
		Addr <=  "0101011000010";
		Trees_din <= x"ff8d2bd5";
		wait for Clk_period;
		Addr <=  "0101011000011";
		Trees_din <= x"6d005708";
		wait for Clk_period;
		Addr <=  "0101011000100";
		Trees_din <= x"de002604";
		wait for Clk_period;
		Addr <=  "0101011000101";
		Trees_din <= x"00502bd5";
		wait for Clk_period;
		Addr <=  "0101011000110";
		Trees_din <= x"00122bd5";
		wait for Clk_period;
		Addr <=  "0101011000111";
		Trees_din <= x"86ff6804";
		wait for Clk_period;
		Addr <=  "0101011001000";
		Trees_din <= x"ffcb2bd5";
		wait for Clk_period;
		Addr <=  "0101011001001";
		Trees_din <= x"00302bd5";
		wait for Clk_period;
		Addr <=  "0101011001010";
		Trees_din <= x"7dffb72c";
		wait for Clk_period;
		Addr <=  "0101011001011";
		Trees_din <= x"4effcc18";
		wait for Clk_period;
		Addr <=  "0101011001100";
		Trees_din <= x"9e000310";
		wait for Clk_period;
		Addr <=  "0101011001101";
		Trees_din <= x"2cff2b08";
		wait for Clk_period;
		Addr <=  "0101011001110";
		Trees_din <= x"00ff4e04";
		wait for Clk_period;
		Addr <=  "0101011001111";
		Trees_din <= x"ffa72bd5";
		wait for Clk_period;
		Addr <=  "0101011010000";
		Trees_din <= x"00482bd5";
		wait for Clk_period;
		Addr <=  "0101011010001";
		Trees_din <= x"c1fe0c04";
		wait for Clk_period;
		Addr <=  "0101011010010";
		Trees_din <= x"00542bd5";
		wait for Clk_period;
		Addr <=  "0101011010011";
		Trees_din <= x"ff932bd5";
		wait for Clk_period;
		Addr <=  "0101011010100";
		Trees_din <= x"dfff8c04";
		wait for Clk_period;
		Addr <=  "0101011010101";
		Trees_din <= x"ffc92bd5";
		wait for Clk_period;
		Addr <=  "0101011010110";
		Trees_din <= x"00762bd5";
		wait for Clk_period;
		Addr <=  "0101011010111";
		Trees_din <= x"0aff9004";
		wait for Clk_period;
		Addr <=  "0101011011000";
		Trees_din <= x"00842bd5";
		wait for Clk_period;
		Addr <=  "0101011011001";
		Trees_din <= x"bbff1608";
		wait for Clk_period;
		Addr <=  "0101011011010";
		Trees_din <= x"dfff9c04";
		wait for Clk_period;
		Addr <=  "0101011011011";
		Trees_din <= x"006c2bd5";
		wait for Clk_period;
		Addr <=  "0101011011100";
		Trees_din <= x"ffe42bd5";
		wait for Clk_period;
		Addr <=  "0101011011101";
		Trees_din <= x"69ff2804";
		wait for Clk_period;
		Addr <=  "0101011011110";
		Trees_din <= x"00092bd5";
		wait for Clk_period;
		Addr <=  "0101011011111";
		Trees_din <= x"ff8d2bd5";
		wait for Clk_period;
		Addr <=  "0101011100000";
		Trees_din <= x"dbff6e0c";
		wait for Clk_period;
		Addr <=  "0101011100001";
		Trees_din <= x"9aff3304";
		wait for Clk_period;
		Addr <=  "0101011100010";
		Trees_din <= x"00242bd5";
		wait for Clk_period;
		Addr <=  "0101011100011";
		Trees_din <= x"e0fe9204";
		wait for Clk_period;
		Addr <=  "0101011100100";
		Trees_din <= x"ffe82bd5";
		wait for Clk_period;
		Addr <=  "0101011100101";
		Trees_din <= x"ff782bd5";
		wait for Clk_period;
		Addr <=  "0101011100110";
		Trees_din <= x"3eff7610";
		wait for Clk_period;
		Addr <=  "0101011100111";
		Trees_din <= x"65fee608";
		wait for Clk_period;
		Addr <=  "0101011101000";
		Trees_din <= x"ac002604";
		wait for Clk_period;
		Addr <=  "0101011101001";
		Trees_din <= x"ffd92bd5";
		wait for Clk_period;
		Addr <=  "0101011101010";
		Trees_din <= x"00662bd5";
		wait for Clk_period;
		Addr <=  "0101011101011";
		Trees_din <= x"28fea904";
		wait for Clk_period;
		Addr <=  "0101011101100";
		Trees_din <= x"003e2bd5";
		wait for Clk_period;
		Addr <=  "0101011101101";
		Trees_din <= x"ffd02bd5";
		wait for Clk_period;
		Addr <=  "0101011101110";
		Trees_din <= x"31ff4708";
		wait for Clk_period;
		Addr <=  "0101011101111";
		Trees_din <= x"bbff8004";
		wait for Clk_period;
		Addr <=  "0101011110000";
		Trees_din <= x"ff812bd5";
		wait for Clk_period;
		Addr <=  "0101011110001";
		Trees_din <= x"00132bd5";
		wait for Clk_period;
		Addr <=  "0101011110010";
		Trees_din <= x"8bffb304";
		wait for Clk_period;
		Addr <=  "0101011110011";
		Trees_din <= x"ffa92bd5";
		wait for Clk_period;
		Addr <=  "0101011110100";
		Trees_din <= x"00482bd5";
		wait for Clk_period;
		Addr <=  "0101011110101";
		Trees_din <= x"1f011f5c";
		wait for Clk_period;
		Addr <=  "0101011110110";
		Trees_din <= x"ab008e28";
		wait for Clk_period;
		Addr <=  "0101011110111";
		Trees_din <= x"7afef808";
		wait for Clk_period;
		Addr <=  "0101011111000";
		Trees_din <= x"b4fe4604";
		wait for Clk_period;
		Addr <=  "0101011111001";
		Trees_din <= x"001c2cb1";
		wait for Clk_period;
		Addr <=  "0101011111010";
		Trees_din <= x"ff7e2cb1";
		wait for Clk_period;
		Addr <=  "0101011111011";
		Trees_din <= x"99ff1210";
		wait for Clk_period;
		Addr <=  "0101011111100";
		Trees_din <= x"20fff708";
		wait for Clk_period;
		Addr <=  "0101011111101";
		Trees_din <= x"5ffead04";
		wait for Clk_period;
		Addr <=  "0101011111110";
		Trees_din <= x"002d2cb1";
		wait for Clk_period;
		Addr <=  "0101011111111";
		Trees_din <= x"ffb82cb1";
		wait for Clk_period;
		Addr <=  "0101100000000";
		Trees_din <= x"31ffb104";
		wait for Clk_period;
		Addr <=  "0101100000001";
		Trees_din <= x"00442cb1";
		wait for Clk_period;
		Addr <=  "0101100000010";
		Trees_din <= x"ffeb2cb1";
		wait for Clk_period;
		Addr <=  "0101100000011";
		Trees_din <= x"c1ff2508";
		wait for Clk_period;
		Addr <=  "0101100000100";
		Trees_din <= x"81ff3c04";
		wait for Clk_period;
		Addr <=  "0101100000101";
		Trees_din <= x"ffbe2cb1";
		wait for Clk_period;
		Addr <=  "0101100000110";
		Trees_din <= x"00292cb1";
		wait for Clk_period;
		Addr <=  "0101100000111";
		Trees_din <= x"aefe8c04";
		wait for Clk_period;
		Addr <=  "0101100001000";
		Trees_din <= x"00382cb1";
		wait for Clk_period;
		Addr <=  "0101100001001";
		Trees_din <= x"ff922cb1";
		wait for Clk_period;
		Addr <=  "0101100001010";
		Trees_din <= x"9dff4a18";
		wait for Clk_period;
		Addr <=  "0101100001011";
		Trees_din <= x"d000da0c";
		wait for Clk_period;
		Addr <=  "0101100001100";
		Trees_din <= x"fcfee208";
		wait for Clk_period;
		Addr <=  "0101100001101";
		Trees_din <= x"28ff4e04";
		wait for Clk_period;
		Addr <=  "0101100001110";
		Trees_din <= x"ffd32cb1";
		wait for Clk_period;
		Addr <=  "0101100001111";
		Trees_din <= x"005b2cb1";
		wait for Clk_period;
		Addr <=  "0101100010000";
		Trees_din <= x"ff7a2cb1";
		wait for Clk_period;
		Addr <=  "0101100010001";
		Trees_din <= x"ac005208";
		wait for Clk_period;
		Addr <=  "0101100010010";
		Trees_din <= x"beffd904";
		wait for Clk_period;
		Addr <=  "0101100010011";
		Trees_din <= x"fffd2cb1";
		wait for Clk_period;
		Addr <=  "0101100010100";
		Trees_din <= x"00712cb1";
		wait for Clk_period;
		Addr <=  "0101100010101";
		Trees_din <= x"ffbb2cb1";
		wait for Clk_period;
		Addr <=  "0101100010110";
		Trees_din <= x"cb005e10";
		wait for Clk_period;
		Addr <=  "0101100010111";
		Trees_din <= x"68fe4908";
		wait for Clk_period;
		Addr <=  "0101100011000";
		Trees_din <= x"1afe7404";
		wait for Clk_period;
		Addr <=  "0101100011001";
		Trees_din <= x"00632cb1";
		wait for Clk_period;
		Addr <=  "0101100011010";
		Trees_din <= x"ff932cb1";
		wait for Clk_period;
		Addr <=  "0101100011011";
		Trees_din <= x"70fee804";
		wait for Clk_period;
		Addr <=  "0101100011100";
		Trees_din <= x"00062cb1";
		wait for Clk_period;
		Addr <=  "0101100011101";
		Trees_din <= x"003f2cb1";
		wait for Clk_period;
		Addr <=  "0101100011110";
		Trees_din <= x"ebfe5b04";
		wait for Clk_period;
		Addr <=  "0101100011111";
		Trees_din <= x"00482cb1";
		wait for Clk_period;
		Addr <=  "0101100100000";
		Trees_din <= x"69fe7104";
		wait for Clk_period;
		Addr <=  "0101100100001";
		Trees_din <= x"00082cb1";
		wait for Clk_period;
		Addr <=  "0101100100010";
		Trees_din <= x"ff7f2cb1";
		wait for Clk_period;
		Addr <=  "0101100100011";
		Trees_din <= x"bdffc50c";
		wait for Clk_period;
		Addr <=  "0101100100100";
		Trees_din <= x"71ffd208";
		wait for Clk_period;
		Addr <=  "0101100100101";
		Trees_din <= x"c2000604";
		wait for Clk_period;
		Addr <=  "0101100100110";
		Trees_din <= x"007d2cb1";
		wait for Clk_period;
		Addr <=  "0101100100111";
		Trees_din <= x"000a2cb1";
		wait for Clk_period;
		Addr <=  "0101100101000";
		Trees_din <= x"fff02cb1";
		wait for Clk_period;
		Addr <=  "0101100101001";
		Trees_din <= x"a2ffca04";
		wait for Clk_period;
		Addr <=  "0101100101010";
		Trees_din <= x"ffa42cb1";
		wait for Clk_period;
		Addr <=  "0101100101011";
		Trees_din <= x"00342cb1";
		wait for Clk_period;
		Addr <=  "0101100101100";
		Trees_din <= x"b1ff0850";
		wait for Clk_period;
		Addr <=  "0101100101101";
		Trees_din <= x"b0ffcf34";
		wait for Clk_period;
		Addr <=  "0101100101110";
		Trees_din <= x"faffa51c";
		wait for Clk_period;
		Addr <=  "0101100101111";
		Trees_din <= x"a3ff020c";
		wait for Clk_period;
		Addr <=  "0101100110000";
		Trees_din <= x"ec001604";
		wait for Clk_period;
		Addr <=  "0101100110001";
		Trees_din <= x"ff8d2dfd";
		wait for Clk_period;
		Addr <=  "0101100110010";
		Trees_din <= x"03ffa904";
		wait for Clk_period;
		Addr <=  "0101100110011";
		Trees_din <= x"ffc82dfd";
		wait for Clk_period;
		Addr <=  "0101100110100";
		Trees_din <= x"00462dfd";
		wait for Clk_period;
		Addr <=  "0101100110101";
		Trees_din <= x"53ff3208";
		wait for Clk_period;
		Addr <=  "0101100110110";
		Trees_din <= x"76ff9d04";
		wait for Clk_period;
		Addr <=  "0101100110111";
		Trees_din <= x"ffcc2dfd";
		wait for Clk_period;
		Addr <=  "0101100111000";
		Trees_din <= x"00612dfd";
		wait for Clk_period;
		Addr <=  "0101100111001";
		Trees_din <= x"43ff7f04";
		wait for Clk_period;
		Addr <=  "0101100111010";
		Trees_din <= x"00222dfd";
		wait for Clk_period;
		Addr <=  "0101100111011";
		Trees_din <= x"ffd52dfd";
		wait for Clk_period;
		Addr <=  "0101100111100";
		Trees_din <= x"e8fec908";
		wait for Clk_period;
		Addr <=  "0101100111101";
		Trees_din <= x"34ffeb04";
		wait for Clk_period;
		Addr <=  "0101100111110";
		Trees_din <= x"00792dfd";
		wait for Clk_period;
		Addr <=  "0101100111111";
		Trees_din <= x"000a2dfd";
		wait for Clk_period;
		Addr <=  "0101101000000";
		Trees_din <= x"d2fe8f08";
		wait for Clk_period;
		Addr <=  "0101101000001";
		Trees_din <= x"6bfee704";
		wait for Clk_period;
		Addr <=  "0101101000010";
		Trees_din <= x"ffb82dfd";
		wait for Clk_period;
		Addr <=  "0101101000011";
		Trees_din <= x"00492dfd";
		wait for Clk_period;
		Addr <=  "0101101000100";
		Trees_din <= x"deff5004";
		wait for Clk_period;
		Addr <=  "0101101000101";
		Trees_din <= x"001c2dfd";
		wait for Clk_period;
		Addr <=  "0101101000110";
		Trees_din <= x"ff8b2dfd";
		wait for Clk_period;
		Addr <=  "0101101000111";
		Trees_din <= x"eaff590c";
		wait for Clk_period;
		Addr <=  "0101101001000";
		Trees_din <= x"2cff2f04";
		wait for Clk_period;
		Addr <=  "0101101001001";
		Trees_din <= x"003d2dfd";
		wait for Clk_period;
		Addr <=  "0101101001010";
		Trees_din <= x"9d000a04";
		wait for Clk_period;
		Addr <=  "0101101001011";
		Trees_din <= x"ff972dfd";
		wait for Clk_period;
		Addr <=  "0101101001100";
		Trees_din <= x"000f2dfd";
		wait for Clk_period;
		Addr <=  "0101101001101";
		Trees_din <= x"0bff7a04";
		wait for Clk_period;
		Addr <=  "0101101001110";
		Trees_din <= x"ffae2dfd";
		wait for Clk_period;
		Addr <=  "0101101001111";
		Trees_din <= x"d1ff0504";
		wait for Clk_period;
		Addr <=  "0101101010000";
		Trees_din <= x"ffc52dfd";
		wait for Clk_period;
		Addr <=  "0101101010001";
		Trees_din <= x"adff1f04";
		wait for Clk_period;
		Addr <=  "0101101010010";
		Trees_din <= x"ffe22dfd";
		wait for Clk_period;
		Addr <=  "0101101010011";
		Trees_din <= x"007e2dfd";
		wait for Clk_period;
		Addr <=  "0101101010100";
		Trees_din <= x"01fe7530";
		wait for Clk_period;
		Addr <=  "0101101010101";
		Trees_din <= x"4dfe5214";
		wait for Clk_period;
		Addr <=  "0101101010110";
		Trees_din <= x"e6000b0c";
		wait for Clk_period;
		Addr <=  "0101101010111";
		Trees_din <= x"8bffc704";
		wait for Clk_period;
		Addr <=  "0101101011000";
		Trees_din <= x"ffcb2dfd";
		wait for Clk_period;
		Addr <=  "0101101011001";
		Trees_din <= x"21ff6704";
		wait for Clk_period;
		Addr <=  "0101101011010";
		Trees_din <= x"fff12dfd";
		wait for Clk_period;
		Addr <=  "0101101011011";
		Trees_din <= x"00722dfd";
		wait for Clk_period;
		Addr <=  "0101101011100";
		Trees_din <= x"36ff5e04";
		wait for Clk_period;
		Addr <=  "0101101011101";
		Trees_din <= x"fff82dfd";
		wait for Clk_period;
		Addr <=  "0101101011110";
		Trees_din <= x"ffad2dfd";
		wait for Clk_period;
		Addr <=  "0101101011111";
		Trees_din <= x"75ffa50c";
		wait for Clk_period;
		Addr <=  "0101101100000";
		Trees_din <= x"79ff2b04";
		wait for Clk_period;
		Addr <=  "0101101100001";
		Trees_din <= x"ffeb2dfd";
		wait for Clk_period;
		Addr <=  "0101101100010";
		Trees_din <= x"9bff5b04";
		wait for Clk_period;
		Addr <=  "0101101100011";
		Trees_din <= x"00822dfd";
		wait for Clk_period;
		Addr <=  "0101101100100";
		Trees_din <= x"00072dfd";
		wait for Clk_period;
		Addr <=  "0101101100101";
		Trees_din <= x"a0ff5708";
		wait for Clk_period;
		Addr <=  "0101101100110";
		Trees_din <= x"21ff9904";
		wait for Clk_period;
		Addr <=  "0101101100111";
		Trees_din <= x"ffec2dfd";
		wait for Clk_period;
		Addr <=  "0101101101000";
		Trees_din <= x"ff9a2dfd";
		wait for Clk_period;
		Addr <=  "0101101101001";
		Trees_din <= x"89000404";
		wait for Clk_period;
		Addr <=  "0101101101010";
		Trees_din <= x"00592dfd";
		wait for Clk_period;
		Addr <=  "0101101101011";
		Trees_din <= x"ffd92dfd";
		wait for Clk_period;
		Addr <=  "0101101101100";
		Trees_din <= x"b3ff7118";
		wait for Clk_period;
		Addr <=  "0101101101101";
		Trees_din <= x"67005310";
		wait for Clk_period;
		Addr <=  "0101101101110";
		Trees_din <= x"86ffa608";
		wait for Clk_period;
		Addr <=  "0101101101111";
		Trees_din <= x"6aff8f04";
		wait for Clk_period;
		Addr <=  "0101101110000";
		Trees_din <= x"ffe62dfd";
		wait for Clk_period;
		Addr <=  "0101101110001";
		Trees_din <= x"ff9a2dfd";
		wait for Clk_period;
		Addr <=  "0101101110010";
		Trees_din <= x"ebff2004";
		wait for Clk_period;
		Addr <=  "0101101110011";
		Trees_din <= x"00402dfd";
		wait for Clk_period;
		Addr <=  "0101101110100";
		Trees_din <= x"ffc32dfd";
		wait for Clk_period;
		Addr <=  "0101101110101";
		Trees_din <= x"a3ffb804";
		wait for Clk_period;
		Addr <=  "0101101110110";
		Trees_din <= x"00072dfd";
		wait for Clk_period;
		Addr <=  "0101101110111";
		Trees_din <= x"00742dfd";
		wait for Clk_period;
		Addr <=  "0101101111000";
		Trees_din <= x"eaff3e04";
		wait for Clk_period;
		Addr <=  "0101101111001";
		Trees_din <= x"ff8d2dfd";
		wait for Clk_period;
		Addr <=  "0101101111010";
		Trees_din <= x"d1ff7d08";
		wait for Clk_period;
		Addr <=  "0101101111011";
		Trees_din <= x"8c000404";
		wait for Clk_period;
		Addr <=  "0101101111100";
		Trees_din <= x"00132dfd";
		wait for Clk_period;
		Addr <=  "0101101111101";
		Trees_din <= x"007a2dfd";
		wait for Clk_period;
		Addr <=  "0101101111110";
		Trees_din <= x"ffa92dfd";
		wait for Clk_period;
		Addr <=  "0101101111111";
		Trees_din <= x"e7ff7b58";
		wait for Clk_period;
		Addr <=  "0101110000000";
		Trees_din <= x"20ff6824";
		wait for Clk_period;
		Addr <=  "0101110000001";
		Trees_din <= x"de00401c";
		wait for Clk_period;
		Addr <=  "0101110000010";
		Trees_din <= x"bbff220c";
		wait for Clk_period;
		Addr <=  "0101110000011";
		Trees_din <= x"1aff0908";
		wait for Clk_period;
		Addr <=  "0101110000100";
		Trees_din <= x"6bfe9904";
		wait for Clk_period;
		Addr <=  "0101110000101";
		Trees_din <= x"ffd42f59";
		wait for Clk_period;
		Addr <=  "0101110000110";
		Trees_din <= x"00652f59";
		wait for Clk_period;
		Addr <=  "0101110000111";
		Trees_din <= x"ffbe2f59";
		wait for Clk_period;
		Addr <=  "0101110001000";
		Trees_din <= x"5cff9108";
		wait for Clk_period;
		Addr <=  "0101110001001";
		Trees_din <= x"49ffa604";
		wait for Clk_period;
		Addr <=  "0101110001010";
		Trees_din <= x"00612f59";
		wait for Clk_period;
		Addr <=  "0101110001011";
		Trees_din <= x"ffe02f59";
		wait for Clk_period;
		Addr <=  "0101110001100";
		Trees_din <= x"b1febe04";
		wait for Clk_period;
		Addr <=  "0101110001101";
		Trees_din <= x"00182f59";
		wait for Clk_period;
		Addr <=  "0101110001110";
		Trees_din <= x"ff852f59";
		wait for Clk_period;
		Addr <=  "0101110001111";
		Trees_din <= x"e9fe2a04";
		wait for Clk_period;
		Addr <=  "0101110010000";
		Trees_din <= x"001e2f59";
		wait for Clk_period;
		Addr <=  "0101110010001";
		Trees_din <= x"ff802f59";
		wait for Clk_period;
		Addr <=  "0101110010010";
		Trees_din <= x"c9ffb714";
		wait for Clk_period;
		Addr <=  "0101110010011";
		Trees_din <= x"00ff0c04";
		wait for Clk_period;
		Addr <=  "0101110010100";
		Trees_din <= x"ff8a2f59";
		wait for Clk_period;
		Addr <=  "0101110010101";
		Trees_din <= x"61ffcc08";
		wait for Clk_period;
		Addr <=  "0101110010110";
		Trees_din <= x"eaff3504";
		wait for Clk_period;
		Addr <=  "0101110010111";
		Trees_din <= x"ffa82f59";
		wait for Clk_period;
		Addr <=  "0101110011000";
		Trees_din <= x"00302f59";
		wait for Clk_period;
		Addr <=  "0101110011001";
		Trees_din <= x"8bffae04";
		wait for Clk_period;
		Addr <=  "0101110011010";
		Trees_din <= x"001e2f59";
		wait for Clk_period;
		Addr <=  "0101110011011";
		Trees_din <= x"ff932f59";
		wait for Clk_period;
		Addr <=  "0101110011100";
		Trees_din <= x"55ffea10";
		wait for Clk_period;
		Addr <=  "0101110011101";
		Trees_din <= x"be002908";
		wait for Clk_period;
		Addr <=  "0101110011110";
		Trees_din <= x"61ffa004";
		wait for Clk_period;
		Addr <=  "0101110011111";
		Trees_din <= x"003c2f59";
		wait for Clk_period;
		Addr <=  "0101110100000";
		Trees_din <= x"ffbf2f59";
		wait for Clk_period;
		Addr <=  "0101110100001";
		Trees_din <= x"03007604";
		wait for Clk_period;
		Addr <=  "0101110100010";
		Trees_din <= x"ff912f59";
		wait for Clk_period;
		Addr <=  "0101110100011";
		Trees_din <= x"00172f59";
		wait for Clk_period;
		Addr <=  "0101110100100";
		Trees_din <= x"17ffd708";
		wait for Clk_period;
		Addr <=  "0101110100101";
		Trees_din <= x"cafe2004";
		wait for Clk_period;
		Addr <=  "0101110100110";
		Trees_din <= x"ffb22f59";
		wait for Clk_period;
		Addr <=  "0101110100111";
		Trees_din <= x"00292f59";
		wait for Clk_period;
		Addr <=  "0101110101000";
		Trees_din <= x"86ffc504";
		wait for Clk_period;
		Addr <=  "0101110101001";
		Trees_din <= x"00642f59";
		wait for Clk_period;
		Addr <=  "0101110101010";
		Trees_din <= x"fff52f59";
		wait for Clk_period;
		Addr <=  "0101110101011";
		Trees_din <= x"7dffb730";
		wait for Clk_period;
		Addr <=  "0101110101100";
		Trees_din <= x"4effcc20";
		wait for Clk_period;
		Addr <=  "0101110101101";
		Trees_din <= x"f9ff0d10";
		wait for Clk_period;
		Addr <=  "0101110101110";
		Trees_din <= x"faff4708";
		wait for Clk_period;
		Addr <=  "0101110101111";
		Trees_din <= x"faff2304";
		wait for Clk_period;
		Addr <=  "0101110110000";
		Trees_din <= x"ffda2f59";
		wait for Clk_period;
		Addr <=  "0101110110001";
		Trees_din <= x"00682f59";
		wait for Clk_period;
		Addr <=  "0101110110010";
		Trees_din <= x"3effb604";
		wait for Clk_period;
		Addr <=  "0101110110011";
		Trees_din <= x"ff9b2f59";
		wait for Clk_period;
		Addr <=  "0101110110100";
		Trees_din <= x"003e2f59";
		wait for Clk_period;
		Addr <=  "0101110110101";
		Trees_din <= x"c1fe4008";
		wait for Clk_period;
		Addr <=  "0101110110110";
		Trees_din <= x"6ffee404";
		wait for Clk_period;
		Addr <=  "0101110110111";
		Trees_din <= x"00612f59";
		wait for Clk_period;
		Addr <=  "0101110111000";
		Trees_din <= x"ffde2f59";
		wait for Clk_period;
		Addr <=  "0101110111001";
		Trees_din <= x"fb003104";
		wait for Clk_period;
		Addr <=  "0101110111010";
		Trees_din <= x"ff882f59";
		wait for Clk_period;
		Addr <=  "0101110111011";
		Trees_din <= x"00002f59";
		wait for Clk_period;
		Addr <=  "0101110111100";
		Trees_din <= x"bbff990c";
		wait for Clk_period;
		Addr <=  "0101110111101";
		Trees_din <= x"0400a608";
		wait for Clk_period;
		Addr <=  "0101110111110";
		Trees_din <= x"01ff0a04";
		wait for Clk_period;
		Addr <=  "0101110111111";
		Trees_din <= x"006e2f59";
		wait for Clk_period;
		Addr <=  "0101111000000";
		Trees_din <= x"ffec2f59";
		wait for Clk_period;
		Addr <=  "0101111000001";
		Trees_din <= x"ffc12f59";
		wait for Clk_period;
		Addr <=  "0101111000010";
		Trees_din <= x"ffb72f59";
		wait for Clk_period;
		Addr <=  "0101111000011";
		Trees_din <= x"dbff6e0c";
		wait for Clk_period;
		Addr <=  "0101111000100";
		Trees_din <= x"9aff3304";
		wait for Clk_period;
		Addr <=  "0101111000101";
		Trees_din <= x"00242f59";
		wait for Clk_period;
		Addr <=  "0101111000110";
		Trees_din <= x"9eff0c04";
		wait for Clk_period;
		Addr <=  "0101111000111";
		Trees_din <= x"ffe02f59";
		wait for Clk_period;
		Addr <=  "0101111001000";
		Trees_din <= x"ff7f2f59";
		wait for Clk_period;
		Addr <=  "0101111001001";
		Trees_din <= x"7f000e10";
		wait for Clk_period;
		Addr <=  "0101111001010";
		Trees_din <= x"65fee608";
		wait for Clk_period;
		Addr <=  "0101111001011";
		Trees_din <= x"2fff2104";
		wait for Clk_period;
		Addr <=  "0101111001100";
		Trees_din <= x"ffaa2f59";
		wait for Clk_period;
		Addr <=  "0101111001101";
		Trees_din <= x"00522f59";
		wait for Clk_period;
		Addr <=  "0101111001110";
		Trees_din <= x"a5ff6904";
		wait for Clk_period;
		Addr <=  "0101111001111";
		Trees_din <= x"000e2f59";
		wait for Clk_period;
		Addr <=  "0101111010000";
		Trees_din <= x"ff9a2f59";
		wait for Clk_period;
		Addr <=  "0101111010001";
		Trees_din <= x"73ffae04";
		wait for Clk_period;
		Addr <=  "0101111010010";
		Trees_din <= x"00252f59";
		wait for Clk_period;
		Addr <=  "0101111010011";
		Trees_din <= x"2eff6604";
		wait for Clk_period;
		Addr <=  "0101111010100";
		Trees_din <= x"ffdf2f59";
		wait for Clk_period;
		Addr <=  "0101111010101";
		Trees_din <= x"ff7c2f59";
		wait for Clk_period;
		Addr <=  "0101111010110";
		Trees_din <= x"01fe7b50";
		wait for Clk_period;
		Addr <=  "0101111010111";
		Trees_din <= x"2cff1f18";
		wait for Clk_period;
		Addr <=  "0101111011000";
		Trees_din <= x"3aff1508";
		wait for Clk_period;
		Addr <=  "0101111011001";
		Trees_din <= x"d6008304";
		wait for Clk_period;
		Addr <=  "0101111011010";
		Trees_din <= x"ff8530b5";
		wait for Clk_period;
		Addr <=  "0101111011011";
		Trees_din <= x"ffe130b5";
		wait for Clk_period;
		Addr <=  "0101111011100";
		Trees_din <= x"70feb408";
		wait for Clk_period;
		Addr <=  "0101111011101";
		Trees_din <= x"67ff4d04";
		wait for Clk_period;
		Addr <=  "0101111011110";
		Trees_din <= x"006430b5";
		wait for Clk_period;
		Addr <=  "0101111011111";
		Trees_din <= x"000830b5";
		wait for Clk_period;
		Addr <=  "0101111100000";
		Trees_din <= x"1fff8904";
		wait for Clk_period;
		Addr <=  "0101111100001";
		Trees_din <= x"fff630b5";
		wait for Clk_period;
		Addr <=  "0101111100010";
		Trees_din <= x"ffa730b5";
		wait for Clk_period;
		Addr <=  "0101111100011";
		Trees_din <= x"b5ff031c";
		wait for Clk_period;
		Addr <=  "0101111100100";
		Trees_din <= x"00ffa20c";
		wait for Clk_period;
		Addr <=  "0101111100101";
		Trees_din <= x"3fffc604";
		wait for Clk_period;
		Addr <=  "0101111100110";
		Trees_din <= x"ff8f30b5";
		wait for Clk_period;
		Addr <=  "0101111100111";
		Trees_din <= x"94ff4204";
		wait for Clk_period;
		Addr <=  "0101111101000";
		Trees_din <= x"003530b5";
		wait for Clk_period;
		Addr <=  "0101111101001";
		Trees_din <= x"ffe830b5";
		wait for Clk_period;
		Addr <=  "0101111101010";
		Trees_din <= x"43ffa908";
		wait for Clk_period;
		Addr <=  "0101111101011";
		Trees_din <= x"7dff9404";
		wait for Clk_period;
		Addr <=  "0101111101100";
		Trees_din <= x"ffd430b5";
		wait for Clk_period;
		Addr <=  "0101111101101";
		Trees_din <= x"005130b5";
		wait for Clk_period;
		Addr <=  "0101111101110";
		Trees_din <= x"1f004804";
		wait for Clk_period;
		Addr <=  "0101111101111";
		Trees_din <= x"ffa130b5";
		wait for Clk_period;
		Addr <=  "0101111110000";
		Trees_din <= x"001a30b5";
		wait for Clk_period;
		Addr <=  "0101111110001";
		Trees_din <= x"9bff6f10";
		wait for Clk_period;
		Addr <=  "0101111110010";
		Trees_din <= x"36fefb08";
		wait for Clk_period;
		Addr <=  "0101111110011";
		Trees_din <= x"47008904";
		wait for Clk_period;
		Addr <=  "0101111110100";
		Trees_din <= x"ffbe30b5";
		wait for Clk_period;
		Addr <=  "0101111110101";
		Trees_din <= x"002930b5";
		wait for Clk_period;
		Addr <=  "0101111110110";
		Trees_din <= x"70fe5d04";
		wait for Clk_period;
		Addr <=  "0101111110111";
		Trees_din <= x"fffc30b5";
		wait for Clk_period;
		Addr <=  "0101111111000";
		Trees_din <= x"006f30b5";
		wait for Clk_period;
		Addr <=  "0101111111001";
		Trees_din <= x"84ffb508";
		wait for Clk_period;
		Addr <=  "0101111111010";
		Trees_din <= x"f5000e04";
		wait for Clk_period;
		Addr <=  "0101111111011";
		Trees_din <= x"005430b5";
		wait for Clk_period;
		Addr <=  "0101111111100";
		Trees_din <= x"ffd430b5";
		wait for Clk_period;
		Addr <=  "0101111111101";
		Trees_din <= x"ff9f30b5";
		wait for Clk_period;
		Addr <=  "0101111111110";
		Trees_din <= x"fbff8b28";
		wait for Clk_period;
		Addr <=  "0101111111111";
		Trees_din <= x"b6ff0b14";
		wait for Clk_period;
		Addr <=  "0110000000000";
		Trees_din <= x"84006a10";
		wait for Clk_period;
		Addr <=  "0110000000001";
		Trees_din <= x"c5ff0308";
		wait for Clk_period;
		Addr <=  "0110000000010";
		Trees_din <= x"9bff3104";
		wait for Clk_period;
		Addr <=  "0110000000011";
		Trees_din <= x"005730b5";
		wait for Clk_period;
		Addr <=  "0110000000100";
		Trees_din <= x"ffcb30b5";
		wait for Clk_period;
		Addr <=  "0110000000101";
		Trees_din <= x"69fee104";
		wait for Clk_period;
		Addr <=  "0110000000110";
		Trees_din <= x"000530b5";
		wait for Clk_period;
		Addr <=  "0110000000111";
		Trees_din <= x"ff7a30b5";
		wait for Clk_period;
		Addr <=  "0110000001000";
		Trees_din <= x"006030b5";
		wait for Clk_period;
		Addr <=  "0110000001001";
		Trees_din <= x"7aff0204";
		wait for Clk_period;
		Addr <=  "0110000001010";
		Trees_din <= x"ffa430b5";
		wait for Clk_period;
		Addr <=  "0110000001011";
		Trees_din <= x"0500a408";
		wait for Clk_period;
		Addr <=  "0110000001100";
		Trees_din <= x"33fee504";
		wait for Clk_period;
		Addr <=  "0110000001101";
		Trees_din <= x"ffd330b5";
		wait for Clk_period;
		Addr <=  "0110000001110";
		Trees_din <= x"003830b5";
		wait for Clk_period;
		Addr <=  "0110000001111";
		Trees_din <= x"5e002f04";
		wait for Clk_period;
		Addr <=  "0110000010000";
		Trees_din <= x"ffb230b5";
		wait for Clk_period;
		Addr <=  "0110000010001";
		Trees_din <= x"003c30b5";
		wait for Clk_period;
		Addr <=  "0110000010010";
		Trees_din <= x"59ffdf20";
		wait for Clk_period;
		Addr <=  "0110000010011";
		Trees_din <= x"41fef310";
		wait for Clk_period;
		Addr <=  "0110000010100";
		Trees_din <= x"5effb608";
		wait for Clk_period;
		Addr <=  "0110000010101";
		Trees_din <= x"88002004";
		wait for Clk_period;
		Addr <=  "0110000010110";
		Trees_din <= x"002e30b5";
		wait for Clk_period;
		Addr <=  "0110000010111";
		Trees_din <= x"ffb330b5";
		wait for Clk_period;
		Addr <=  "0110000011000";
		Trees_din <= x"65ffaa04";
		wait for Clk_period;
		Addr <=  "0110000011001";
		Trees_din <= x"ff8330b5";
		wait for Clk_period;
		Addr <=  "0110000011010";
		Trees_din <= x"fff230b5";
		wait for Clk_period;
		Addr <=  "0110000011011";
		Trees_din <= x"88000708";
		wait for Clk_period;
		Addr <=  "0110000011100";
		Trees_din <= x"2cffc604";
		wait for Clk_period;
		Addr <=  "0110000011101";
		Trees_din <= x"ffb530b5";
		wait for Clk_period;
		Addr <=  "0110000011110";
		Trees_din <= x"001c30b5";
		wait for Clk_period;
		Addr <=  "0110000011111";
		Trees_din <= x"49ffda04";
		wait for Clk_period;
		Addr <=  "0110000100000";
		Trees_din <= x"ffd030b5";
		wait for Clk_period;
		Addr <=  "0110000100001";
		Trees_din <= x"005830b5";
		wait for Clk_period;
		Addr <=  "0110000100010";
		Trees_din <= x"62ff2610";
		wait for Clk_period;
		Addr <=  "0110000100011";
		Trees_din <= x"15ff3908";
		wait for Clk_period;
		Addr <=  "0110000100100";
		Trees_din <= x"d9ffe604";
		wait for Clk_period;
		Addr <=  "0110000100101";
		Trees_din <= x"ffef30b5";
		wait for Clk_period;
		Addr <=  "0110000100110";
		Trees_din <= x"006e30b5";
		wait for Clk_period;
		Addr <=  "0110000100111";
		Trees_din <= x"70fe5d04";
		wait for Clk_period;
		Addr <=  "0110000101000";
		Trees_din <= x"002530b5";
		wait for Clk_period;
		Addr <=  "0110000101001";
		Trees_din <= x"ff9630b5";
		wait for Clk_period;
		Addr <=  "0110000101010";
		Trees_din <= x"1f006b04";
		wait for Clk_period;
		Addr <=  "0110000101011";
		Trees_din <= x"ff7230b5";
		wait for Clk_period;
		Addr <=  "0110000101100";
		Trees_din <= x"fff230b5";
		wait for Clk_period;
		Addr <=  "0110000101101";
		Trees_din <= x"bbfff964";
		wait for Clk_period;
		Addr <=  "0110000101110";
		Trees_din <= x"1aff3538";
		wait for Clk_period;
		Addr <=  "0110000101111";
		Trees_din <= x"2efff01c";
		wait for Clk_period;
		Addr <=  "0110000110000";
		Trees_din <= x"49ff720c";
		wait for Clk_period;
		Addr <=  "0110000110001";
		Trees_din <= x"71ff9c08";
		wait for Clk_period;
		Addr <=  "0110000110010";
		Trees_din <= x"4eff2704";
		wait for Clk_period;
		Addr <=  "0110000110011";
		Trees_din <= x"ffdb31a1";
		wait for Clk_period;
		Addr <=  "0110000110100";
		Trees_din <= x"005b31a1";
		wait for Clk_period;
		Addr <=  "0110000110101";
		Trees_din <= x"ffa731a1";
		wait for Clk_period;
		Addr <=  "0110000110110";
		Trees_din <= x"88ff9508";
		wait for Clk_period;
		Addr <=  "0110000110111";
		Trees_din <= x"19feec04";
		wait for Clk_period;
		Addr <=  "0110000111000";
		Trees_din <= x"002e31a1";
		wait for Clk_period;
		Addr <=  "0110000111001";
		Trees_din <= x"ff9e31a1";
		wait for Clk_period;
		Addr <=  "0110000111010";
		Trees_din <= x"bcff6d04";
		wait for Clk_period;
		Addr <=  "0110000111011";
		Trees_din <= x"000b31a1";
		wait for Clk_period;
		Addr <=  "0110000111100";
		Trees_din <= x"ffd931a1";
		wait for Clk_period;
		Addr <=  "0110000111101";
		Trees_din <= x"6bfe720c";
		wait for Clk_period;
		Addr <=  "0110000111110";
		Trees_din <= x"71ff9008";
		wait for Clk_period;
		Addr <=  "0110000111111";
		Trees_din <= x"6cfed104";
		wait for Clk_period;
		Addr <=  "0110001000000";
		Trees_din <= x"000131a1";
		wait for Clk_period;
		Addr <=  "0110001000001";
		Trees_din <= x"ff8a31a1";
		wait for Clk_period;
		Addr <=  "0110001000010";
		Trees_din <= x"003d31a1";
		wait for Clk_period;
		Addr <=  "0110001000011";
		Trees_din <= x"83ff2308";
		wait for Clk_period;
		Addr <=  "0110001000100";
		Trees_din <= x"b1ff4304";
		wait for Clk_period;
		Addr <=  "0110001000101";
		Trees_din <= x"001931a1";
		wait for Clk_period;
		Addr <=  "0110001000110";
		Trees_din <= x"ff9931a1";
		wait for Clk_period;
		Addr <=  "0110001000111";
		Trees_din <= x"06ff0a04";
		wait for Clk_period;
		Addr <=  "0110001001000";
		Trees_din <= x"ffee31a1";
		wait for Clk_period;
		Addr <=  "0110001001001";
		Trees_din <= x"005931a1";
		wait for Clk_period;
		Addr <=  "0110001001010";
		Trees_din <= x"9aff570c";
		wait for Clk_period;
		Addr <=  "0110001001011";
		Trees_din <= x"cdffd404";
		wait for Clk_period;
		Addr <=  "0110001001100";
		Trees_din <= x"ffc531a1";
		wait for Clk_period;
		Addr <=  "0110001001101";
		Trees_din <= x"20ffb204";
		wait for Clk_period;
		Addr <=  "0110001001110";
		Trees_din <= x"001a31a1";
		wait for Clk_period;
		Addr <=  "0110001001111";
		Trees_din <= x"007931a1";
		wait for Clk_period;
		Addr <=  "0110001010000";
		Trees_din <= x"0bffce10";
		wait for Clk_period;
		Addr <=  "0110001010001";
		Trees_din <= x"b7004108";
		wait for Clk_period;
		Addr <=  "0110001010010";
		Trees_din <= x"a0ff7a04";
		wait for Clk_period;
		Addr <=  "0110001010011";
		Trees_din <= x"ff7631a1";
		wait for Clk_period;
		Addr <=  "0110001010100";
		Trees_din <= x"fff631a1";
		wait for Clk_period;
		Addr <=  "0110001010101";
		Trees_din <= x"2cff4004";
		wait for Clk_period;
		Addr <=  "0110001010110";
		Trees_din <= x"005a31a1";
		wait for Clk_period;
		Addr <=  "0110001010111";
		Trees_din <= x"ffc931a1";
		wait for Clk_period;
		Addr <=  "0110001011000";
		Trees_din <= x"43ff9808";
		wait for Clk_period;
		Addr <=  "0110001011001";
		Trees_din <= x"39fff704";
		wait for Clk_period;
		Addr <=  "0110001011010";
		Trees_din <= x"003b31a1";
		wait for Clk_period;
		Addr <=  "0110001011011";
		Trees_din <= x"ff9c31a1";
		wait for Clk_period;
		Addr <=  "0110001011100";
		Trees_din <= x"a0ff7d04";
		wait for Clk_period;
		Addr <=  "0110001011101";
		Trees_din <= x"ff8a31a1";
		wait for Clk_period;
		Addr <=  "0110001011110";
		Trees_din <= x"000731a1";
		wait for Clk_period;
		Addr <=  "0110001011111";
		Trees_din <= x"01fe7810";
		wait for Clk_period;
		Addr <=  "0110001100000";
		Trees_din <= x"d8003508";
		wait for Clk_period;
		Addr <=  "0110001100001";
		Trees_din <= x"76fffb04";
		wait for Clk_period;
		Addr <=  "0110001100010";
		Trees_din <= x"fffa31a1";
		wait for Clk_period;
		Addr <=  "0110001100011";
		Trees_din <= x"005a31a1";
		wait for Clk_period;
		Addr <=  "0110001100100";
		Trees_din <= x"1eff5604";
		wait for Clk_period;
		Addr <=  "0110001100101";
		Trees_din <= x"ffee31a1";
		wait for Clk_period;
		Addr <=  "0110001100110";
		Trees_din <= x"ffab31a1";
		wait for Clk_period;
		Addr <=  "0110001100111";
		Trees_din <= x"ff8c31a1";
		wait for Clk_period;
		Addr <=  "0110001101000";
		Trees_din <= x"ab011358";
		wait for Clk_period;
		Addr <=  "0110001101001";
		Trees_din <= x"fcfebc1c";
		wait for Clk_period;
		Addr <=  "0110001101010";
		Trees_din <= x"65ff5e14";
		wait for Clk_period;
		Addr <=  "0110001101011";
		Trees_din <= x"dcff7d08";
		wait for Clk_period;
		Addr <=  "0110001101100";
		Trees_din <= x"cdffd204";
		wait for Clk_period;
		Addr <=  "0110001101101";
		Trees_din <= x"ffda32a5";
		wait for Clk_period;
		Addr <=  "0110001101110";
		Trees_din <= x"006032a5";
		wait for Clk_period;
		Addr <=  "0110001101111";
		Trees_din <= x"dc006f08";
		wait for Clk_period;
		Addr <=  "0110001110000";
		Trees_din <= x"0a008404";
		wait for Clk_period;
		Addr <=  "0110001110001";
		Trees_din <= x"ff8232a5";
		wait for Clk_period;
		Addr <=  "0110001110010";
		Trees_din <= x"fffd32a5";
		wait for Clk_period;
		Addr <=  "0110001110011";
		Trees_din <= x"002932a5";
		wait for Clk_period;
		Addr <=  "0110001110100";
		Trees_din <= x"86ff9a04";
		wait for Clk_period;
		Addr <=  "0110001110101";
		Trees_din <= x"ff8132a5";
		wait for Clk_period;
		Addr <=  "0110001110110";
		Trees_din <= x"ffe332a5";
		wait for Clk_period;
		Addr <=  "0110001110111";
		Trees_din <= x"b1ff141c";
		wait for Clk_period;
		Addr <=  "0110001111000";
		Trees_din <= x"a8002310";
		wait for Clk_period;
		Addr <=  "0110001111001";
		Trees_din <= x"f8ffd508";
		wait for Clk_period;
		Addr <=  "0110001111010";
		Trees_din <= x"effed104";
		wait for Clk_period;
		Addr <=  "0110001111011";
		Trees_din <= x"004132a5";
		wait for Clk_period;
		Addr <=  "0110001111100";
		Trees_din <= x"ff8a32a5";
		wait for Clk_period;
		Addr <=  "0110001111101";
		Trees_din <= x"53ff3404";
		wait for Clk_period;
		Addr <=  "0110001111110";
		Trees_din <= x"003932a5";
		wait for Clk_period;
		Addr <=  "0110001111111";
		Trees_din <= x"000132a5";
		wait for Clk_period;
		Addr <=  "0110010000000";
		Trees_din <= x"eaff5b04";
		wait for Clk_period;
		Addr <=  "0110010000001";
		Trees_din <= x"ffcd32a5";
		wait for Clk_period;
		Addr <=  "0110010000010";
		Trees_din <= x"3eff6504";
		wait for Clk_period;
		Addr <=  "0110010000011";
		Trees_din <= x"000b32a5";
		wait for Clk_period;
		Addr <=  "0110010000100";
		Trees_din <= x"008b32a5";
		wait for Clk_period;
		Addr <=  "0110010000101";
		Trees_din <= x"6d002410";
		wait for Clk_period;
		Addr <=  "0110010000110";
		Trees_din <= x"cfff9c08";
		wait for Clk_period;
		Addr <=  "0110010000111";
		Trees_din <= x"defff204";
		wait for Clk_period;
		Addr <=  "0110010001000";
		Trees_din <= x"005732a5";
		wait for Clk_period;
		Addr <=  "0110010001001";
		Trees_din <= x"ffbd32a5";
		wait for Clk_period;
		Addr <=  "0110010001010";
		Trees_din <= x"76fff504";
		wait for Clk_period;
		Addr <=  "0110010001011";
		Trees_din <= x"ffa932a5";
		wait for Clk_period;
		Addr <=  "0110010001100";
		Trees_din <= x"fffc32a5";
		wait for Clk_period;
		Addr <=  "0110010001101";
		Trees_din <= x"4f003f08";
		wait for Clk_period;
		Addr <=  "0110010001110";
		Trees_din <= x"9dffe104";
		wait for Clk_period;
		Addr <=  "0110010001111";
		Trees_din <= x"fffd32a5";
		wait for Clk_period;
		Addr <=  "0110010010000";
		Trees_din <= x"003d32a5";
		wait for Clk_period;
		Addr <=  "0110010010001";
		Trees_din <= x"8fff8a04";
		wait for Clk_period;
		Addr <=  "0110010010010";
		Trees_din <= x"ff9932a5";
		wait for Clk_period;
		Addr <=  "0110010010011";
		Trees_din <= x"002132a5";
		wait for Clk_period;
		Addr <=  "0110010010100";
		Trees_din <= x"73000018";
		wait for Clk_period;
		Addr <=  "0110010010101";
		Trees_din <= x"64ff0f10";
		wait for Clk_period;
		Addr <=  "0110010010110";
		Trees_din <= x"11ff9108";
		wait for Clk_period;
		Addr <=  "0110010010111";
		Trees_din <= x"41ff4004";
		wait for Clk_period;
		Addr <=  "0110010011000";
		Trees_din <= x"ffae32a5";
		wait for Clk_period;
		Addr <=  "0110010011001";
		Trees_din <= x"002232a5";
		wait for Clk_period;
		Addr <=  "0110010011010";
		Trees_din <= x"afffb904";
		wait for Clk_period;
		Addr <=  "0110010011011";
		Trees_din <= x"007332a5";
		wait for Clk_period;
		Addr <=  "0110010011100";
		Trees_din <= x"000c32a5";
		wait for Clk_period;
		Addr <=  "0110010011101";
		Trees_din <= x"6e009504";
		wait for Clk_period;
		Addr <=  "0110010011110";
		Trees_din <= x"ff8932a5";
		wait for Clk_period;
		Addr <=  "0110010011111";
		Trees_din <= x"000732a5";
		wait for Clk_period;
		Addr <=  "0110010100000";
		Trees_din <= x"ceff4f04";
		wait for Clk_period;
		Addr <=  "0110010100001";
		Trees_din <= x"ffd732a5";
		wait for Clk_period;
		Addr <=  "0110010100010";
		Trees_din <= x"baff8204";
		wait for Clk_period;
		Addr <=  "0110010100011";
		Trees_din <= x"fff432a5";
		wait for Clk_period;
		Addr <=  "0110010100100";
		Trees_din <= x"37ff3d04";
		wait for Clk_period;
		Addr <=  "0110010100101";
		Trees_din <= x"fff032a5";
		wait for Clk_period;
		Addr <=  "0110010100110";
		Trees_din <= x"f1ff4d04";
		wait for Clk_period;
		Addr <=  "0110010100111";
		Trees_din <= x"002632a5";
		wait for Clk_period;
		Addr <=  "0110010101000";
		Trees_din <= x"008b32a5";
		wait for Clk_period;
		Addr <=  "0110010101001";
		Trees_din <= x"89008270";
		wait for Clk_period;
		Addr <=  "0110010101010";
		Trees_din <= x"03ff6430";
		wait for Clk_period;
		Addr <=  "0110010101011";
		Trees_din <= x"0dff9018";
		wait for Clk_period;
		Addr <=  "0110010101100";
		Trees_din <= x"d5ffc808";
		wait for Clk_period;
		Addr <=  "0110010101101";
		Trees_din <= x"fafedc04";
		wait for Clk_period;
		Addr <=  "0110010101110";
		Trees_din <= x"002133f1";
		wait for Clk_period;
		Addr <=  "0110010101111";
		Trees_din <= x"ff8d33f1";
		wait for Clk_period;
		Addr <=  "0110010110000";
		Trees_din <= x"e0ff4a08";
		wait for Clk_period;
		Addr <=  "0110010110001";
		Trees_din <= x"44004604";
		wait for Clk_period;
		Addr <=  "0110010110010";
		Trees_din <= x"004033f1";
		wait for Clk_period;
		Addr <=  "0110010110011";
		Trees_din <= x"ffbc33f1";
		wait for Clk_period;
		Addr <=  "0110010110100";
		Trees_din <= x"13001904";
		wait for Clk_period;
		Addr <=  "0110010110101";
		Trees_din <= x"003a33f1";
		wait for Clk_period;
		Addr <=  "0110010110110";
		Trees_din <= x"ffb733f1";
		wait for Clk_period;
		Addr <=  "0110010110111";
		Trees_din <= x"6a000210";
		wait for Clk_period;
		Addr <=  "0110010111000";
		Trees_din <= x"98ff8208";
		wait for Clk_period;
		Addr <=  "0110010111001";
		Trees_din <= x"1afe5804";
		wait for Clk_period;
		Addr <=  "0110010111010";
		Trees_din <= x"ffe233f1";
		wait for Clk_period;
		Addr <=  "0110010111011";
		Trees_din <= x"ff7233f1";
		wait for Clk_period;
		Addr <=  "0110010111100";
		Trees_din <= x"1eff3904";
		wait for Clk_period;
		Addr <=  "0110010111101";
		Trees_din <= x"006a33f1";
		wait for Clk_period;
		Addr <=  "0110010111110";
		Trees_din <= x"ffaa33f1";
		wait for Clk_period;
		Addr <=  "0110010111111";
		Trees_din <= x"8bffd404";
		wait for Clk_period;
		Addr <=  "0110011000000";
		Trees_din <= x"005633f1";
		wait for Clk_period;
		Addr <=  "0110011000001";
		Trees_din <= x"ffd633f1";
		wait for Clk_period;
		Addr <=  "0110011000010";
		Trees_din <= x"82ff7820";
		wait for Clk_period;
		Addr <=  "0110011000011";
		Trees_din <= x"b4feea10";
		wait for Clk_period;
		Addr <=  "0110011000100";
		Trees_din <= x"0efe8e08";
		wait for Clk_period;
		Addr <=  "0110011000101";
		Trees_din <= x"8dfdc204";
		wait for Clk_period;
		Addr <=  "0110011000110";
		Trees_din <= x"ffb833f1";
		wait for Clk_period;
		Addr <=  "0110011000111";
		Trees_din <= x"004e33f1";
		wait for Clk_period;
		Addr <=  "0110011001000";
		Trees_din <= x"64fefa04";
		wait for Clk_period;
		Addr <=  "0110011001001";
		Trees_din <= x"003033f1";
		wait for Clk_period;
		Addr <=  "0110011001010";
		Trees_din <= x"ffd133f1";
		wait for Clk_period;
		Addr <=  "0110011001011";
		Trees_din <= x"9aff6208";
		wait for Clk_period;
		Addr <=  "0110011001100";
		Trees_din <= x"a4ff5504";
		wait for Clk_period;
		Addr <=  "0110011001101";
		Trees_din <= x"005a33f1";
		wait for Clk_period;
		Addr <=  "0110011001110";
		Trees_din <= x"ffd433f1";
		wait for Clk_period;
		Addr <=  "0110011001111";
		Trees_din <= x"6dffed04";
		wait for Clk_period;
		Addr <=  "0110011010000";
		Trees_din <= x"ff9533f1";
		wait for Clk_period;
		Addr <=  "0110011010001";
		Trees_din <= x"ffde33f1";
		wait for Clk_period;
		Addr <=  "0110011010010";
		Trees_din <= x"20ff8e10";
		wait for Clk_period;
		Addr <=  "0110011010011";
		Trees_din <= x"2fff2508";
		wait for Clk_period;
		Addr <=  "0110011010100";
		Trees_din <= x"01fed604";
		wait for Clk_period;
		Addr <=  "0110011010101";
		Trees_din <= x"ff9a33f1";
		wait for Clk_period;
		Addr <=  "0110011010110";
		Trees_din <= x"003433f1";
		wait for Clk_period;
		Addr <=  "0110011010111";
		Trees_din <= x"9affb704";
		wait for Clk_period;
		Addr <=  "0110011011000";
		Trees_din <= x"fffe33f1";
		wait for Clk_period;
		Addr <=  "0110011011001";
		Trees_din <= x"006f33f1";
		wait for Clk_period;
		Addr <=  "0110011011010";
		Trees_din <= x"33ffbd08";
		wait for Clk_period;
		Addr <=  "0110011011011";
		Trees_din <= x"42ff7e04";
		wait for Clk_period;
		Addr <=  "0110011011100";
		Trees_din <= x"ffb433f1";
		wait for Clk_period;
		Addr <=  "0110011011101";
		Trees_din <= x"000d33f1";
		wait for Clk_period;
		Addr <=  "0110011011110";
		Trees_din <= x"6fff7f04";
		wait for Clk_period;
		Addr <=  "0110011011111";
		Trees_din <= x"006b33f1";
		wait for Clk_period;
		Addr <=  "0110011100000";
		Trees_din <= x"ffe833f1";
		wait for Clk_period;
		Addr <=  "0110011100001";
		Trees_din <= x"02fea718";
		wait for Clk_period;
		Addr <=  "0110011100010";
		Trees_din <= x"a8ff8f10";
		wait for Clk_period;
		Addr <=  "0110011100011";
		Trees_din <= x"2a01260c";
		wait for Clk_period;
		Addr <=  "0110011100100";
		Trees_din <= x"faffcc08";
		wait for Clk_period;
		Addr <=  "0110011100101";
		Trees_din <= x"cdff4f04";
		wait for Clk_period;
		Addr <=  "0110011100110";
		Trees_din <= x"fffc33f1";
		wait for Clk_period;
		Addr <=  "0110011100111";
		Trees_din <= x"007b33f1";
		wait for Clk_period;
		Addr <=  "0110011101000";
		Trees_din <= x"ffec33f1";
		wait for Clk_period;
		Addr <=  "0110011101001";
		Trees_din <= x"ffdc33f1";
		wait for Clk_period;
		Addr <=  "0110011101010";
		Trees_din <= x"2fff9104";
		wait for Clk_period;
		Addr <=  "0110011101011";
		Trees_din <= x"ffb233f1";
		wait for Clk_period;
		Addr <=  "0110011101100";
		Trees_din <= x"003033f1";
		wait for Clk_period;
		Addr <=  "0110011101101";
		Trees_din <= x"29ffa510";
		wait for Clk_period;
		Addr <=  "0110011101110";
		Trees_din <= x"4dfdec04";
		wait for Clk_period;
		Addr <=  "0110011101111";
		Trees_din <= x"003833f1";
		wait for Clk_period;
		Addr <=  "0110011110000";
		Trees_din <= x"34004908";
		wait for Clk_period;
		Addr <=  "0110011110001";
		Trees_din <= x"8800ff04";
		wait for Clk_period;
		Addr <=  "0110011110010";
		Trees_din <= x"ff7f33f1";
		wait for Clk_period;
		Addr <=  "0110011110011";
		Trees_din <= x"001933f1";
		wait for Clk_period;
		Addr <=  "0110011110100";
		Trees_din <= x"002833f1";
		wait for Clk_period;
		Addr <=  "0110011110101";
		Trees_din <= x"e9feaf04";
		wait for Clk_period;
		Addr <=  "0110011110110";
		Trees_din <= x"ffd733f1";
		wait for Clk_period;
		Addr <=  "0110011110111";
		Trees_din <= x"42ff3904";
		wait for Clk_period;
		Addr <=  "0110011111000";
		Trees_din <= x"ffe433f1";
		wait for Clk_period;
		Addr <=  "0110011111001";
		Trees_din <= x"beffb404";
		wait for Clk_period;
		Addr <=  "0110011111010";
		Trees_din <= x"001833f1";
		wait for Clk_period;
		Addr <=  "0110011111011";
		Trees_din <= x"007833f1";
		wait for Clk_period;
		Addr <=  "0110011111100";
		Trees_din <= x"0000001f";
		wait for Clk_period;

        -- Reset valid flag
        Valid_node <= '0';
        wait for Clk_period; 
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101010000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111000000101";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111001101101";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "0000000101101110";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "0000000011100001";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111010011000";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111000010000";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111001010000";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111010100100";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111001111111";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111010110011";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111001111100";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "0000000101000001";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111001101011";
        wait for Clk_period; 
        Features_din <= "0000000011111111";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111110111101111";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111001001000";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111000001010";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111001101001";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111010010111";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111001101101";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "0000001000011000";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111010110011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111010011111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111110110010110";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111001111001";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111010001110";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "0000000010111110";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "1111110111101010";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111010100100";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111000111111";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111001001010";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111110111110101";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111110111011000";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111010100101";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "0000000110100101";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111000101101";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110110100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111001010011";
        wait for Clk_period; 
        Features_din <= "1111111010101110";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "0000000011000110";
        wait for Clk_period; 
        Features_din <= "0000000011100001";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "0000000011100001";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111000011010";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111111001011000";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "0000000011011000";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "0000000011010101";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111001000010";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111001100101";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "0000000011111001";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "1111111001100111";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111001000000";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111010001011";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111001111101";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "0000000100000000";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111010010001";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111010001110";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111001101011";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111001001001";
        wait for Clk_period; 
        Features_din <= "1111111001110101";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111010011001";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111001101111";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000010111100";
        wait for Clk_period; 
        Features_din <= "0000000101011011";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111000111011";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111001101000";
        wait for Clk_period; 
        Features_din <= "1111111000101000";
        wait for Clk_period; 
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111001100011";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "0000001011011000";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "1111111001100100";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(6, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000000101010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "0000000011101000";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111001100110";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111010000111";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "0000000100010100";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "0000000011000000";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111010001111";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111010010101";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "0000000011000000";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111000110001";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111010101110";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "0000000011010111";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111000011101";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000011101100";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "0000000100111001";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111110111100100";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(5, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101100001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111001011001";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "1111111010011001";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111010011000";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111010011011";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "0000000100100011";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111001111011";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111010001110";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111001100000";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111000111011";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111010110011";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111110111011011";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "1111111010000001";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "1111111001111110";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111000001101";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "0000000011111111";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111001010000";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111000110110";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111001101010";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111001101100";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000000011100101";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111010011000";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "0000000011000001";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111001101010";
        wait for Clk_period; 
        Features_din <= "1111111000000010";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "0000001011011110";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111100110010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111010000001";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "0000000100100111";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111001010101";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111010000110";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "0000000011100110";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111010010111";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111001010001";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111001110001";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111000110000";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "0000000010111000";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111001001010";
        wait for Clk_period; 
        Features_din <= "1111111000111101";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "0000001001011001";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111010011000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111100111001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111000111111";
        wait for Clk_period; 
        Features_din <= "1111111010001101";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "0000000011100110";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111010100101";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111001111011";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "0000000010111101";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111010100101";
        wait for Clk_period; 
        Features_din <= "1111111001101001";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "0000000011011000";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111001101001";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111010000100";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111010001110";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111010011011";
        wait for Clk_period; 
        Features_din <= "1111111001010011";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111001001101";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111000110001";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111010110011";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "0000001010100101";
        wait for Clk_period; 
        Features_din <= "1111111000110101";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(5, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000000001000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111001110101";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "0000000011000001";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111000000110";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111010101000";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111001011111";
        wait for Clk_period; 
        Features_din <= "0000000011110010";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111010001011";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111001001111";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "0000000011111100";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111001001001";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111000111101";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111000101110";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111010000100";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111001010111";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111110111111000";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111000100101";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "0000000011000000";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "1111111000001010";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111010100101";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "0000001011010100";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101000101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111001010000";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111001011101";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111001100110";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111010000001";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111001011100";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111001011000";
        wait for Clk_period; 
        Features_din <= "1111111010011010";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111010001100";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111001111011";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111010001011";
        wait for Clk_period; 
        Features_din <= "1111111010101010";
        wait for Clk_period; 
        Features_din <= "0000000100101000";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000011110011";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "1111111001111101";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "0000000100001100";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111110111110101";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111001001100";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111001110001";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111010011111";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111000111010";
        wait for Clk_period; 
        Features_din <= "1111111001110111";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000011100011";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111001100001";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111001100011";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111000110010";
        wait for Clk_period; 
        Features_din <= "1111111000001100";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "0000001001000111";
        wait for Clk_period; 
        Features_din <= "1111111010010101";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000000001011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "0000000010111110";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111110111100001";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111110110001101";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111110101111000";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "0000000100101110";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111000101001";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111001010100";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111000110001";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "0000000100000011";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111010000011";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "1111111001101111";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "0000000101101011";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111010011010";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111010010101";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111001111000";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "1111110111111110";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111010000110";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "0000001000011001";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101111101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "1111111000101111";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "0000000100001000";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111010101000";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "0000000011011100";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111010001111";
        wait for Clk_period; 
        Features_din <= "1111110111000110";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111010011111";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111001011101";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111010010011";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111001110111";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111010011110";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111000111010";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111001111001";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "0000000010111000";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111001011011";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111001100111";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111001001001";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "0000001011101011";
        wait for Clk_period; 
        Features_din <= "1111111001011000";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111100111010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111110111110111";
        wait for Clk_period; 
        Features_din <= "0000000010101100";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111001110000";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111010001011";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "0000000011011000";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111010100100";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111010010000";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111010010000";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111010001010";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111010011000";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111000001010";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111010100100";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "1111111000000001";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111001000010";
        wait for Clk_period; 
        Features_din <= "1111111010101000";
        wait for Clk_period; 
        Features_din <= "1111111001011100";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111010000001";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000011010101";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111010101000";
        wait for Clk_period; 
        Features_din <= "0000000010101100";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "0000000011000001";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111000110101";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111000111000";
        wait for Clk_period; 
        Features_din <= "1111111010010101";
        wait for Clk_period; 
        Features_din <= "1111111001000010";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "0000001001000000";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000000010011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010000100";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "1111111010010011";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111111000101100";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111000000000";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "0000000011000100";
        wait for Clk_period; 
        Features_din <= "0000000011111010";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "0000000011110111";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111000111000";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111111010011110";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "0000000100011111";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111000001101";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "0000000011000010";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111010000001";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "0000000011001100";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111010001010";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111000111111";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111010100000";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111010010111";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "0000000011000000";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010111101";
        wait for Clk_period; 
        Features_din <= "0000000010101101";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "0000000011101010";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111001110101";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "0000000010110010";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "0000001001001111";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110111000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "0000000011101010";
        wait for Clk_period; 
        Features_din <= "0000000011010101";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "0000000011111001";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111000000010";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "0000000100001001";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111000101010";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111010010111";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111010011110";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111001011110";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111001100111";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111001010011";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111110100000110";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "0000000010111101";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111010100000";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111000011010";
        wait for Clk_period; 
        Features_din <= "1111111010011011";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111010010101";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111110111001110";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111010100000";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "0000000110111001";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111001010000";
        wait for Clk_period; 
        Features_din <= "1111111000000101";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "0000001011100110";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101100001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010010001";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "0000000100001000";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111110111100100";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "0000000100011010";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111000110111";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "0000000110011100";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111010101110";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111010110011";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111010100101";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111001001001";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111010000011";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "0000000011001100";
        wait for Clk_period; 
        Features_din <= "0000000011011011";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111110110101111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111001111110";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111001010010";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111010011111";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111010100101";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111001110000";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111001000100";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111010011111";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "0000000011010111";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111010001010";
        wait for Clk_period; 
        Features_din <= "1111111001010111";
        wait for Clk_period; 
        Features_din <= "1111111010011010";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "0000001011111100";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111100000011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "0000000101010111";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "0000000101111011";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111010101110";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111001100011";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "0000000011010101";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111001100101";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111000111000";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111010000000";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111000110010";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111001011011";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111010001101";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111110111101111";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111010001110";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111001110011";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "0000000100001101";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111010011111";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111010000111";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111001010101";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "0000000011010001";
        wait for Clk_period; 
        Features_din <= "0000000011111100";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111110111001111";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111010001111";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111001101101";
        wait for Clk_period; 
        Features_din <= "1111111001101111";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "0000000111111011";
        wait for Clk_period; 
        Features_din <= "1111111000110010";
        wait for Clk_period; 
        Features_din <= "1111111010001110";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110110000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111000101100";
        wait for Clk_period; 
        Features_din <= "1111111001011000";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "0000000100100011";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "0000000011101101";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111001000100";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111010011000";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111000010110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "0000000100011010";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111010101000";
        wait for Clk_period; 
        Features_din <= "1111110111110101";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111001100101";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111000100101";
        wait for Clk_period; 
        Features_din <= "1111111010010111";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111000100000";
        wait for Clk_period; 
        Features_din <= "1111111001100100";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111001110100";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111001110111";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111000011011";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111010011110";
        wait for Clk_period; 
        Features_din <= "1111111000101111";
        wait for Clk_period; 
        Features_din <= "1111111001011011";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "0000001001010000";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110010110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111000010101";
        wait for Clk_period; 
        Features_din <= "1111111010011000";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "0000000100101100";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "1111111001011100";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "1111111001011111";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111001001001";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "0000000011101101";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111111010100000";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111010000111";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "0000000011101100";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111001111001";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111001011110";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "0000000010111101";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000100100101";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111000000011";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111001001111";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111010010011";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000100000101";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "0000000011001111";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "0000000011001011";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111010000111";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "0000001011001001";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110100000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111000011101";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "0000000110011110";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111001101110";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111010010000";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111010110011";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111010011000";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111010000110";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "0000000011000100";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111001000000";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111010000010";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "0000000011011011";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111110101110011";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "0000000100100101";
        wait for Clk_period; 
        Features_din <= "0000000011111010";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000010111100";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "0000001000110000";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111001011110";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111000100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111000010010";
        wait for Clk_period; 
        Features_din <= "1111111001100000";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "0000000011101110";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "1111111010011110";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111001001101";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111111000001100";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111010000010";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111010000011";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "0000000011001010";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111010001101";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "1111110111111001";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111010101000";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111010000111";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111010010011";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "0000000100011110";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "1111111000010000";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111001101000";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "0000000010110010";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111010000000";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "0000000011001101";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111010000010";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111000101010";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111000011000";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111000111101";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111001010010";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "1111111010011111";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111001110101";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111010011010";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "1111111001111010";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111001111101";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "0000000011111101";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111001111110";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111001111101";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "0000001000110101";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111010001111";
        wait for Clk_period; 
        Features_din <= "0000000011000000";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101110101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111001111011";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "0000000011110111";
        wait for Clk_period; 
        Features_din <= "0000000011001110";
        wait for Clk_period; 
        Features_din <= "1111110111110110";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111110111110000";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000011011111";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111001101111";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "1111111010001011";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "0000000011000101";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111010011000";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "0000000011111010";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111010001110";
        wait for Clk_period; 
        Features_din <= "1111111001000100";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111110111110111";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111001001101";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "0000000011110100";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111000001010";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111000101010";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111110110000111";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111010001001";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111001101011";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111001111110";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111001000010";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111010001111";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111001001111";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "0000000100010101";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111010001001";
        wait for Clk_period; 
        Features_din <= "1111111001101011";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111001000001";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "0000001001101011";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110000001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111010101110";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "0000000011001100";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "0000000100010110";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "0000000010110011";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111000101101";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000100011000";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111110111110000";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111110111001101";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111010001010";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000100101100";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111000011010";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "0000000011000000";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000011110000";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111001110101";
        wait for Clk_period; 
        Features_din <= "1111111000110101";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "0000001011000000";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111010101110";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110010001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111001111110";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "0000000011000100";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "0000000100100100";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "1111111010000011";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111001110010";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "0000000011101101";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "0000000011001000";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "0000000011101101";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "0000000010110010";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "0000000011011101";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111110110011011";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "0000000010101100";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111010001100";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111001111000";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111010100000";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111001100011";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111001110100";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111001011100";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111001000010";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111010000010";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111010000111";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111000101000";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000100011001";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111001001110";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000100010011";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111001010000";
        wait for Clk_period; 
        Features_din <= "1111111001101101";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "0000001011100110";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "0000000011110010";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101101011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111110111111001";
        wait for Clk_period; 
        Features_din <= "1111111001100110";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111110111101010";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111010000110";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "0000000010101101";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111110111011110";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000011001011";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111001011011";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111000101001";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111110111100111";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111001110001";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111010000110";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "0000000010111101";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111110110101111";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111010010111";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111001110100";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111001011100";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111010000111";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111001001100";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111001100100";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "0000000011000100";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "0000001100000010";
        wait for Clk_period; 
        Features_din <= "1111111010011111";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "0000000011011111";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(6, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110010010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111000000111";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "0000000011110000";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111001110010";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111001111001";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "0000000110000011";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111001100000";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "0000000011001110";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111010000100";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111001101100";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111000101110";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111001101011";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111010011010";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111001011100";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111010001110";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111010010101";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111010001111";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "0000000011010000";
        wait for Clk_period; 
        Features_din <= "0000000010110010";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "1111111000111111";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111001101011";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111000011100";
        wait for Clk_period; 
        Features_din <= "1111111001110111";
        wait for Clk_period; 
        Features_din <= "1111111001111000";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "0000000110010111";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111001101000";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101110100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111001110111";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "0000000011001011";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111001010101";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111001011101";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "0000000100111110";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111000000010";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111010101010";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111010000000";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111110111010111";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "0000000101101000";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111010100101";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111001101100";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111010000010";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111010001101";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "0000000100111010";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000010110011";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111001100101";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111001100111";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111010001001";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "1111111010010101";
        wait for Clk_period; 
        Features_din <= "0000000100001111";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110100100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "0000000011010000";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "0000000100000100";
        wait for Clk_period; 
        Features_din <= "1111111001111011";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111000111001";
        wait for Clk_period; 
        Features_din <= "0000000011101101";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111001101111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "0000000011010110";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111010001101";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111000011011";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111001101110";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111111010011000";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111001011010";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111010011010";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111010001001";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111010010001";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111001010111";
        wait for Clk_period; 
        Features_din <= "1111111001111000";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "0000000011110011";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "1111110111010001";
        wait for Clk_period; 
        Features_din <= "0000000011010110";
        wait for Clk_period; 
        Features_din <= "1111111001001011";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111010010111";
        wait for Clk_period; 
        Features_din <= "1111111010000111";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111010010101";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111010001100";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111000000001";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111000000010";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111010101110";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000010111111";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "0000000100100110";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111010011110";
        wait for Clk_period; 
        Features_din <= "1111111000001101";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "0000001001101011";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "0000000011011000";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111100101011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111010110011";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "1111111010010101";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111001010001";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "1111111001101011";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111001110101";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111010101000";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111010011000";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111000111000";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111001111111";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111001110100";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111000111111";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "0000000011001000";
        wait for Clk_period; 
        Features_din <= "0000000010101100";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111001001000";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111001101001";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111010000100";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "1111111010000111";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "1111111001101010";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111010100000";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "0000000010111111";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "0000000111110100";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110011011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "0000000010110011";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "1111111000101100";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111010101010";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "0000000010101100";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "0000000100100111";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "0000000100000101";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111001110011";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "0000000011111001";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111001010010";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111001110111";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "0000000011101001";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111000011101";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111010010111";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "0000001000010001";
        wait for Clk_period; 
        Features_din <= "1111111001101100";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111010010011";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "1111111010100000";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111101101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111001011010";
        wait for Clk_period; 
        Features_din <= "1111111000011100";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111111001010101";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111001011111";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000000011011011";
        wait for Clk_period; 
        Features_din <= "1111111010000010";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "0000000010101101";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000011000111";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111001111100";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "1111111001110011";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "0000000100010011";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111000010001";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111110110100110";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "1111111010000000";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111000111100";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111010010101";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111001000101";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111001001000";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111001001110";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111001100011";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111001011000";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111001111100";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111010000001";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000010111000";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000011101001";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "0000000100011010";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111000101101";
        wait for Clk_period; 
        Features_din <= "1111111001100110";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "0000001001100110";
        wait for Clk_period; 
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "1111111001110000";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101100110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "0000000100000111";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111000110000";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111010001111";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111000011100";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111010011010";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111010101010";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111001111111";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "0000000011011001";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111111000000000";
        wait for Clk_period; 
        Features_din <= "1111111010000111";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "0000001000110110";
        wait for Clk_period; 
        Features_din <= "1111111010001001";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101100110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111001110000";
        wait for Clk_period; 
        Features_din <= "1111111001010111";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "0000000010101100";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111110111010000";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111000001110";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111010100000";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111000011111";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111000100111";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111010000011";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111001101100";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111010010000";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111001110010";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "0000000011000010";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111010010111";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111001100100";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111000101110";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000001011100110";
        wait for Clk_period; 
        Features_din <= "1111111000100111";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111010000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111100001111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111001010001";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010111101";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111000110100";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000010101101";
        wait for Clk_period; 
        Features_din <= "0000000011000001";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "0000000011001100";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "0000000011001011";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111010110011";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111010001011";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111010010111";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111001110100";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111001101010";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111010000100";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111001001001";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111000111001";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111010011000";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111001110111";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "0000000011110111";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "0000000100010011";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111001101111";
        wait for Clk_period; 
        Features_din <= "1111111010001001";
        wait for Clk_period; 
        Features_din <= "1111111010000110";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "0000001010100010";
        wait for Clk_period; 
        Features_din <= "1111111010001100";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "0000000011000111";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101110111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010010000";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "0000000011101010";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111110110000000";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000101111111";
        wait for Clk_period; 
        Features_din <= "1111111010100100";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111110111010111";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111010011001";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111000100110";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111000101110";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "0000000011001100";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111001101000";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "0000000011100010";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111001110010";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111000101010";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111000111010";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111000110110";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111010100000";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111001101111";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111001111000";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111010000010";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111000100111";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111001111011";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111001111011";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111010000000";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "0000001000111100";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110101111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111010101010";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "0000000011100101";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "0000000011000001";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "0000000010111100";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111010010001";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111001111110";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111001000100";
        wait for Clk_period; 
        Features_din <= "1111111010100000";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "0000000111011101";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "1111111001101111";
        wait for Clk_period; 
        Features_din <= "1111111010000110";
        wait for Clk_period; 
        Features_din <= "1111111010100101";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111010011010";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111110111011111";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111111000111000";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111010100000";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111000110111";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111001110001";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111110110110111";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111010001011";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111010110011";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "0000000010110010";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111001110111";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111001010011";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "1111111001101011";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111001011011";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111010001110";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "0000001000010011";
        wait for Clk_period; 
        Features_din <= "1111111000111101";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(3, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111100101100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111001101101";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "0000000011011011";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "0000000011001001";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111001000101";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111000111011";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "1111111010100101";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000100101111";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111000101011";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111000000011";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111001010101";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111001101111";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "0000000011000000";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111010100000";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111001111101";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "0000000010111000";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111010010001";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "1111111001100110";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111001100100";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111001011111";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111000010001";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000000100001010";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111010010000";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "0000000011010010";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "0000001011111101";
        wait for Clk_period; 
        Features_din <= "1111111010000010";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "0000000011111110";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(6, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110011111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "0000000011000101";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "1111111001111001";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "0000000101010100";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111001000001";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111001100101";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "0000000011000010";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "0000000011000111";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111001011111";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "0000000100001010";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111001100001";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111001000010";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111010010101";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111001001111";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111001010011";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111010010001";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111010010000";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111010011001";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "0000000101101110";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "0000001011101001";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111001011101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000000011101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111000110001";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "0000000010101100";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "0000000011011011";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111001110010";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111001101111";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000010111101";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111001000111";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111001011110";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111010000100";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111010010111";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "0000000011011000";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111001101100";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111001110000";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "0000000011010010";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111001001111";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000011010101";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111010000111";
        wait for Clk_period; 
        Features_din <= "1111111001010000";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111010000011";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111010101110";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111001001110";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111010011000";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111001111000";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "0000001001110001";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101010111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111001111110";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111110111010000";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "0000000100110111";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111000111000";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "0000000010111110";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111001101100";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111001001110";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "0000000011101010";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111000111100";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111010011001";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111010000000";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "0000000100000101";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "0000000011011101";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111000000111";
        wait for Clk_period; 
        Features_din <= "1111111001111110";
        wait for Clk_period; 
        Features_din <= "1111110110010001";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "0000001001100100";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111010000111";
        wait for Clk_period; 
        Features_din <= "0000000011000111";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000011000111";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111010011000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110010010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111001100000";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "0000000011011100";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "1111111010000111";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111010110011";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "0000000011001101";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "0000000011010000";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111010001100";
        wait for Clk_period; 
        Features_din <= "1111111001101001";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "0000000011111100";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111010011001";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111110111101001";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111010101010";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "0000000011010010";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111010000000";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "0000000100111010";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111110111101110";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111001111110";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111010010101";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "0000000011110010";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "0000000011011101";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111000000101";
        wait for Clk_period; 
        Features_din <= "1111111001010101";
        wait for Clk_period; 
        Features_din <= "1111111001001000";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "0000001000011111";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111100010101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "1111111000011001";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111010000100";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111000011110";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "0000000011000111";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111001110111";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111010001111";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111110101000100";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111111010001101";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111010101010";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "0000001000101100";
        wait for Clk_period; 
        Features_din <= "1111111000110011";
        wait for Clk_period; 
        Features_din <= "1111111001111011";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101011001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010000001";
        wait for Clk_period; 
        Features_din <= "1111111010001100";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111001101111";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "0000000010111101";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111001000101";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111110111000100";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "0000000011101010";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111010011011";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111010010011";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111001011100";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111001111111";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111010001001";
        wait for Clk_period; 
        Features_din <= "1111111010011110";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111001110000";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111010011001";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111001010010";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "0000000100000110";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000011000000";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111010011111";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111000011011";
        wait for Clk_period; 
        Features_din <= "1111111010010011";
        wait for Clk_period; 
        Features_din <= "1111111001010111";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "0000001001011101";
        wait for Clk_period; 
        Features_din <= "1111111010011001";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "0000000011000010";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000011101100";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111100110001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "0000000010110011";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111001010110";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000000011001010";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "0000000011010101";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "0000000100000111";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111001110011";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111000100111";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111001110111";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111001101100";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111010010000";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000011001010";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111000100000";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111000010110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111110110110100";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111000011000";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111010001111";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111010000111";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000011011101";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111010010101";
        wait for Clk_period; 
        Features_din <= "1111111001001111";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111000011101";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111010110011";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101001111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111010101110";
        wait for Clk_period; 
        Features_din <= "1111111001011111";
        wait for Clk_period; 
        Features_din <= "0000000011111110";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111001111100";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111010001011";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111001011001";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111110111101110";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111010011111";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111001110011";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111001101000";
        wait for Clk_period; 
        Features_din <= "0000000101010110";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111001111011";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111001111011";
        wait for Clk_period; 
        Features_din <= "0000000011100110";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111001100101";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111010001011";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111110111001100";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111000010110";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111000011010";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111010101000";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111000011100";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111000111110";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111000010100";
        wait for Clk_period; 
        Features_din <= "0000000011000110";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111001100011";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "0000000010110010";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "0000000111110011";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "0000000011100010";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111000110010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101011100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111001111000";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "0000000010111101";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "1111111010001110";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "0000000011000100";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "0000000011011011";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111001110011";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111000010111";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "0000000011001010";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111001101001";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "0000000010111100";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "0000000011011000";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111110111101100";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111001111011";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111001110010";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111010010011";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111010100100";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "1111111010100100";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000011110110";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111010101000";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111001010001";
        wait for Clk_period; 
        Features_din <= "1111111010100101";
        wait for Clk_period; 
        Features_din <= "1111111010010011";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101110110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111010100000";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "0000000011001100";
        wait for Clk_period; 
        Features_din <= "0000000011001010";
        wait for Clk_period; 
        Features_din <= "1111111001111011";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111000010000";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111010100101";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "0000000011011010";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111010100000";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111000100111";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111001111000";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111010101110";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111000100010";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111001000011";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111001101100";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111001000100";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111001011100";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "0000000100110011";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111110111101010";
        wait for Clk_period; 
        Features_din <= "1111111000101110";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111001111111";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "0000000100101000";
        wait for Clk_period; 
        Features_din <= "1111110110011001";
        wait for Clk_period; 
        Features_din <= "1111111000110000";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101011100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "1111111001100110";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "0000000011111100";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111001011000";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111001010101";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "0000000100011011";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111010000011";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111110111101101";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111000111110";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111000101001";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111010100000";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111001111000";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111001100000";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111001000011";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101010011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "0000000100000000";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "0000000101000010";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111010000100";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "0000000101000110";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "0000000010111110";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111001000011";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000011010010";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "0000000011111100";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "0000000010110011";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111010010000";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111010001101";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "0000000011101111";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111001110000";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "1111110111110110";
        wait for Clk_period; 
        Features_din <= "1111111000101111";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "0000000011101111";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "0000000110101100";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111001000100";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "0000000011010101";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111010010000";
        wait for Clk_period; 
        Features_din <= "1111111001111101";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111001111101";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111010100000";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111001111001";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000100101111";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "0000000101101001";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111010001100";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111010001100";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "1111111001110100";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111000010111";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "0000001100011001";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "0000000010110010";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "0000000011010010";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(5, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110111100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111001110001";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "0000000100001010";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111010010011";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111001010010";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111010010001";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "0000000011110101";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "0000000011001110";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "0000000010110011";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "0000000011110100";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111001110010";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111110111011111";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111010001101";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "0000000011100000";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111001010111";
        wait for Clk_period; 
        Features_din <= "1111111001011011";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "1111111001101111";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "0000000111101000";
        wait for Clk_period; 
        Features_din <= "1111111000010110";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111010010111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110001000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "1111110111100110";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "1111111000011011";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111001100110";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "0000000011100100";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111001010110";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111110111010101";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111010000010";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111001011101";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111010001010";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111001111011";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111000000101";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111010011010";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111010011011";
        wait for Clk_period; 
        Features_din <= "1111111001010111";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111010100101";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111010010111";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "1111111010010111";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111001011101";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111001101010";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111001010010";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "0000001011101101";
        wait for Clk_period; 
        Features_din <= "1111111001111001";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000100101000";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110100100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111001110011";
        wait for Clk_period; 
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "0000000100001100";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111000001111";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111000101101";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "0000000100001010";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111010101110";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111010010101";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "0000000100010010";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111000110111";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111001011011";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111001111110";
        wait for Clk_period; 
        Features_din <= "1111111010101010";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111001001000";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111001001011";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111001110001";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111001011110";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111110111010101";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111001011011";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "0000000011010111";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000000100111110";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111010001111";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111001000100";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "1111111001110001";
        wait for Clk_period; 
        Features_din <= "1111111000110000";
        wait for Clk_period; 
        Features_din <= "1111111000111111";
        wait for Clk_period; 
        Features_din <= "1111111001010100";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "0000001100110000";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "0000000100000111";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110001110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111001000001";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "0000000011100001";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "0000000011000010";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "1111111001100111";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111000001000";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111010101010";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000010111000";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111010001001";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111001000000";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111000011101";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111010101000";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111001111000";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111001100000";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111001000111";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000011010001";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111010001001";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111011101100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111110110000001";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "0000000111010010";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111010011001";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111010011001";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111110110100010";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111010001010";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111001101011";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "0000000011101000";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111010001010";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111001110101";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111001100011";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111000110001";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111010001100";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111010001001";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "0000000100011010";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110100010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010001100";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111010010101";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111000100110";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111001100000";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "0000000100000110";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "0000000100110100";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111010001110";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111000010111";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111001110100";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111001001101";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111001100011";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111001011111";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111001001101";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "0000000100011000";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111000100101";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111001001101";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "0000001011101111";
        wait for Clk_period; 
        Features_din <= "1111111001010111";
        wait for Clk_period; 
        Features_din <= "1111111010000100";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000000000001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111010100100";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "0000000100010001";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "0000000011001101";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "1111111010011111";
        wait for Clk_period; 
        Features_din <= "0000000011000010";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111010000111";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111001001001";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111010000000";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111010011000";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111001101100";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111010101010";
        wait for Clk_period; 
        Features_din <= "1111111010011110";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "0000000011010011";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "0000000011001101";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111001100110";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111001100111";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111010010000";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111000100000";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "0000000011010110";
        wait for Clk_period; 
        Features_din <= "0000000101111101";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111000101101";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111010110011";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111010100100";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111001101001";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111001000100";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111010001110";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111010011110";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "0000000011100101";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111001111010";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000000101110001";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111010010011";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111010000011";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111010000100";
        wait for Clk_period; 
        Features_din <= "1111111010001010";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111011010011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111001100000";
        wait for Clk_period; 
        Features_din <= "1111111010101010";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "0000000100101110";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111000101111";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111110110011010";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "0000000011000100";
        wait for Clk_period; 
        Features_din <= "1111111001101110";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111000011111";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111000000001";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000011110111";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111010101010";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111000111110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111001111011";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111001100011";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111001101110";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "0000000011100000";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111010101000";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111110101100101";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111110111011001";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111001110000";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111001110100";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111010010111";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111001000011";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111111001001001";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "0000000100100001";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111001101011";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111010000010";
        wait for Clk_period; 
        Features_din <= "1111111010000001";
        wait for Clk_period; 
        Features_din <= "1111111001000111";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "1111111010011000";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "0000001100010100";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "0000000010111110";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111011001010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000011011011";
        wait for Clk_period; 
        Features_din <= "1111111001000010";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "0000000011000001";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111010100100";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "0000000011100101";
        wait for Clk_period; 
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111001001011";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111010011110";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111010011110";
        wait for Clk_period; 
        Features_din <= "1111111001001000";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111010010001";
        wait for Clk_period; 
        Features_din <= "1111111010000111";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "0000001000100111";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111001101110";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111010010001";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101011001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111110101001110";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "0000000011111010";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111010110011";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111010000011";
        wait for Clk_period; 
        Features_din <= "1111111001110010";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "0000000011110001";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111110111010100";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111010001001";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "0000000100001110";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111010000000";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111010001101";
        wait for Clk_period; 
        Features_din <= "1111111010001111";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111110111101111";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111000111010";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111010110011";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111000110001";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111001110100";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111010010011";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111010011001";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111010000000";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000100100000";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111010011010";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111000100111";
        wait for Clk_period; 
        Features_din <= "1111111010001111";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111000111110";
        wait for Clk_period; 
        Features_din <= "1111111001111111";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111010101110";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "0000000011001010";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111001111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111010001010";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111001111001";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "0000000101011010";
        wait for Clk_period; 
        Features_din <= "1111111000100000";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000011110001";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "0000000101000100";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111001010001";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111001111111";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111010010000";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111001000001";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "0000000011000001";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111001101010";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "0000000011100110";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111010100100";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111010001101";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111001111010";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "0000000011000110";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111000011011";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111010001111";
        wait for Clk_period; 
        Features_din <= "1111111010011110";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111010001101";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000110101101";
        wait for Clk_period; 
        Features_din <= "1111111010000000";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101011100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "0000000011000101";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "1111111001111111";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111010000000";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "1111111001111110";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111010000001";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "0000000011000111";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "0000000011000010";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "0000000110011011";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111001010010";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111000110110";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "0000000100000101";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111010001010";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111110111111101";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000011100011";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111001011001";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111001101100";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111000011001";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111001110000";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111001101101";
        wait for Clk_period; 
        Features_din <= "1111111001011010";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "1111111001001111";
        wait for Clk_period; 
        Features_din <= "1111111010000001";
        wait for Clk_period; 
        Features_din <= "1111111001010011";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "0000001001010000";
        wait for Clk_period; 
        Features_din <= "1111111010011001";
        wait for Clk_period; 
        Features_din <= "1111111001111110";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101101101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "1111111010011000";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "0000000011111111";
        wait for Clk_period; 
        Features_din <= "0000000010111101";
        wait for Clk_period; 
        Features_din <= "1111111001010111";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000010110011";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "0000000011101101";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "0000000101010101";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111110111101110";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111001110111";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111010011111";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111000110011";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111001000011";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111010000100";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111010011110";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111010000110";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111010000000";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111001101111";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000000011101101";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "1111111001111011";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111010011011";
        wait for Clk_period; 
        Features_din <= "1111111001000110";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111110111101101";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111001111101";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "0000000011011001";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "0000001010010001";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111001100100";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111011101010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "0000000011110111";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111001010011";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111001001000";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111010000001";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "0000000100111100";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "0000000011101111";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "0000000011000100";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "1111111010010001";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "0000000100111010";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "0000000011011110";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111001110011";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111001011111";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111111001000011";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111000011011";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111010001011";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111010000110";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111111001000000";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111000111100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000000011001100";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "1111111000110110";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000001001101101";
        wait for Clk_period; 
        Features_din <= "1111111001100101";
        wait for Clk_period; 
        Features_din <= "1111111000101110";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "0000000011101100";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111100101011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111001101011";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "0000000110001000";
        wait for Clk_period; 
        Features_din <= "1111111001000001";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "0000000011111001";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "0000000011010000";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111010100000";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "0000000100000001";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111001110111";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111001101100";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "1111111010011011";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111001111111";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111001110111";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111000101000";
        wait for Clk_period; 
        Features_din <= "1111111001100100";
        wait for Clk_period; 
        Features_din <= "1111111010101010";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111010100100";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "0000001000110111";
        wait for Clk_period; 
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110000011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111001110011";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "0000000011001111";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111000111011";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111001001001";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "1111111001001011";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111001100000";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111001111010";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "1111111010101110";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "0000000011011000";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111000101101";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "0000000101011110";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111000101011";
        wait for Clk_period; 
        Features_din <= "1111111000010110";
        wait for Clk_period; 
        Features_din <= "1111111010001001";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111001111011";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111000000011";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111000110011";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111001011101";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "0000000011001110";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111001000001";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111010011010";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111110110001111";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111000100111";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111001110111";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000011100110";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111001011000";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111010001010";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "1111111010001010";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "0000001001010000";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "0000000011111010";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111011110101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000011001101";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111001110000";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111010010111";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111000111011";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "0000000011001101";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "0000000100000101";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111000011110";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111010101000";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "0000000011100111";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111010011010";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111000111011";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111000000011";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111010010101";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "0000000011001011";
        wait for Clk_period; 
        Features_din <= "1111111000111100";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111001001110";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111001100110";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111001111011";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111001001000";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111001101100";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111001111111";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111001011111";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "0000000110001101";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "0000000011100011";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "0000000011110110";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110111011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111000111011";
        wait for Clk_period; 
        Features_din <= "1111111001110000";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "0000000011110011";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "0000000011001100";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111000110111";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111110110110110";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111010011011";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "0000000011001000";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111001111000";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111001010110";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111001011010";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111110111010000";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111000110001";
        wait for Clk_period; 
        Features_din <= "1111111001110001";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "0000000011100110";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "0000000011100011";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111001000010";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111010011011";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111000011100";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111001001000";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111110110110111";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111001000110";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111111001001100";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111001111111";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111010001110";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111001110010";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "0000000011000100";
        wait for Clk_period; 
        Features_din <= "0000000100110001";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111001100100";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "1111111010000010";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "1111111010100100";
        wait for Clk_period; 
        Features_din <= "1111111001010110";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111010110011";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "0000001000011110";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111011110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "0000000100001101";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "0000000100011011";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111110111111110";
        wait for Clk_period; 
        Features_din <= "0000000011001100";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111110101101000";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111001100110";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "0000000100000100";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111010011000";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "0000000100010110";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111001001101";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "0000000011010011";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111010011011";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111010000011";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111000001101";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111010011111";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111111010000000";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111010011001";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "0000000011011000";
        wait for Clk_period; 
        Features_din <= "0000000100101000";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111001110011";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111010000010";
        wait for Clk_period; 
        Features_din <= "1111111001110111";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111001101111";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111000010100";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000100100001";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "0000000011111000";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "1111111001001011";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111000010100";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "0000001011110010";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101010000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "1111111010010001";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "0000000100001010";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "1111111001111110";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111001001101";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "0000000011000000";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "0000000100010000";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111010100101";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "1111111010010000";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111010000110";
        wait for Clk_period; 
        Features_din <= "1111111001100000";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111010011111";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "0000000011001001";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111110110100110";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111001110000";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111000101111";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000100011010";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000011100000";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111001010000";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000001100010011";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110010011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000011111100";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "0000000011001001";
        wait for Clk_period; 
        Features_din <= "0000000010111110";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111001011111";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111010100101";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111010011111";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111001010111";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "0000000011001011";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111000111001";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111000001101";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "0000000011000101";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111001000001";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111001111100";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111010000110";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111001010001";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111110111101010";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111001000100";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000000100000101";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111001011101";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111001010111";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111110110010111";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "0000001100001101";
        wait for Clk_period; 
        Features_din <= "1111111001011010";
        wait for Clk_period; 
        Features_din <= "1111111010001011";
        wait for Clk_period; 
        Features_din <= "0000000011000100";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "0000000011001110";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101001000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000011001000";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111110100010011";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "0000000110000100";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111001100110";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "0000000011011000";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111001001000";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "0000000011001000";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111001111101";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111001010110";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111111001001010";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111001110010";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111110110101110";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "1111111010010111";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111001101101";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101011101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111000111100";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111001100101";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "0000000011000110";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111010001010";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111000110100";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111000001110";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111001011011";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111001100011";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111001011100";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111001011100";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111001001101";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000000100000100";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111010010111";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "0000000010111000";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "0000000011001010";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111000101001";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111010100000";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000001010111111";
        wait for Clk_period; 
        Features_din <= "1111110111101000";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000000011100110";
        wait for Clk_period; 
        Features_din <= "1111111010000001";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111000101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010001001";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "1111111001100111";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111000001011";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "0000000011011100";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "0000000101000100";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111010010000";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111001111010";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "0000000011110110";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111010011001";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111010101110";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000011110111";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111110110110101";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111001101011";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "0000000011000000";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111010001001";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111010001110";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111010011010";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111001111111";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111000110011";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "0000000011010011";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111001001011";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111001110011";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111001110111";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "0000001011110000";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(3, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111111111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111110111110100";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "0000000101000000";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "0000000101011110";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111010011000";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111110111000100";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111010101010";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111110111010001";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111010110011";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111001001001";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111010000000";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111001110000";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111010000100";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111001011111";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "0000000101100000";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111001111101";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101101000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111001011111";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111010100000";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111010000011";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111010010101";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "0000000100111110";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111001001001";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "0000000100111110";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111001111100";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "0000000011000010";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111010011111";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111010000110";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111010010000";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "1111111010101000";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111010100100";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "1111111010001101";
        wait for Clk_period; 
        Features_din <= "1111111001011010";
        wait for Clk_period; 
        Features_din <= "1111111000111001";
        wait for Clk_period; 
        Features_din <= "1111111001100111";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "0000001001110010";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111100011110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010011011";
        wait for Clk_period; 
        Features_din <= "1111111010000011";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111010110011";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111001001111";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111000111100";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "0000000011101111";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111000101110";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "0000000011011100";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111110111100001";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111010000100";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111000111100";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111001110010";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111001001001";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "0000000100000100";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "1111111001011011";
        wait for Clk_period; 
        Features_din <= "1111110111101100";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111010000011";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "0000001011010110";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101100001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111001111100";
        wait for Clk_period; 
        Features_din <= "1111111001010001";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "0000000100001101";
        wait for Clk_period; 
        Features_din <= "0000000011100111";
        wait for Clk_period; 
        Features_din <= "1111111001000110";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111000101101";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111010100101";
        wait for Clk_period; 
        Features_din <= "0000000011010101";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "0000000011010111";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111001110011";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111010001111";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111000101010";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111110111011000";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111001010000";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111010001011";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111010011111";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "0000000100000111";
        wait for Clk_period; 
        Features_din <= "0000000010110010";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111110111011101";
        wait for Clk_period; 
        Features_din <= "1111111000111000";
        wait for Clk_period; 
        Features_din <= "1111110111111010";
        wait for Clk_period; 
        Features_din <= "1111111000011101";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "0000000111111010";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111001010110";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "0000000010111100";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110110000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010010001";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "0000000011001110";
        wait for Clk_period; 
        Features_din <= "0000000010110011";
        wait for Clk_period; 
        Features_din <= "1111111010001111";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111001000110";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "1111111001101110";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "0000000011011011";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111111001100001";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111010001001";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111001101100";
        wait for Clk_period; 
        Features_din <= "1111111000100100";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111000101110";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111010010001";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111010011001";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111111010110011";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111001101010";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111001101000";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111010001111";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111111010011011";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111010001110";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000011001001";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "0000000011000001";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "0000000100011010";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111001000100";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "0000001011101000";
        wait for Clk_period; 
        Features_din <= "1111111000111111";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111100100100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "0000000011111000";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111010010111";
        wait for Clk_period; 
        Features_din <= "1111111001001011";
        wait for Clk_period; 
        Features_din <= "1111111001110000";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111010011010";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111001100110";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111010101010";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111010000110";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111010000000";
        wait for Clk_period; 
        Features_din <= "1111111010001001";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111010000110";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111010000011";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111000000111";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "0000000010101100";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "0000000011011100";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111000001000";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "0000000011000100";
        wait for Clk_period; 
        Features_din <= "0000000011010101";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "0000000010111100";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111010101010";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111000100000";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111000011101";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111000101010";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111000101011";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111010110011";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "0000001011011001";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "0000000011001010";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110011001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010011000";
        wait for Clk_period; 
        Features_din <= "1111111001001110";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "0000000011101011";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "0000000011001000";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111111010011110";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111000101110";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111001011011";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111001111000";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111001111001";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111010001101";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111010010101";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "0000000100001001";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111110111100000";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111010101000";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "0000000010111110";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111111001111001";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111010100100";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111010011000";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "1111111010000111";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111010000011";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111001100110";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111010011011";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111010010011";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111000101111";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000101011110";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111010001001";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111010000010";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111110111110010";
        wait for Clk_period; 
        Features_din <= "1111110111100000";
        wait for Clk_period; 
        Features_din <= "1111111000011100";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "0000001001110010";
        wait for Clk_period; 
        Features_din <= "1111111000101001";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "0000000010101100";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(5, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110001000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111110111010010";
        wait for Clk_period; 
        Features_din <= "1111111001111001";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "0000000100101111";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "1111111010001100";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111010000011";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111010001101";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "0000000011001110";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111001101001";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "0000000011110011";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111010001010";
        wait for Clk_period; 
        Features_din <= "1111111001011000";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111001001100";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "0000000100001110";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111001111101";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111010101110";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111010010101";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "0000000011000100";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111110101111011";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111010000100";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111001101001";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111001100000";
        wait for Clk_period; 
        Features_din <= "1111111001101100";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111010000000";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111000001100";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111111000101101";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111001101100";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111000111010";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111010101110";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111111010101110";
        wait for Clk_period; 
        Features_din <= "1111111010110011";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "0000001010010011";
        wait for Clk_period; 
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "0000000011000000";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "0000000010110011";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110010101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111001010101";
        wait for Clk_period; 
        Features_din <= "1111111010100101";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "0000000011010111";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "1111111010001101";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111000100000";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111010101010";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111010010011";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "0000000010101100";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "0000000010101100";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "1111111010010001";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "1111111000101111";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111001011011";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111001111100";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111001101100";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000000011010011";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111010010001";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111000111011";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111000101100";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111001011110";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111000101101";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000011110110";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111010011001";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111001110011";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "0000001010101011";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111100111100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111001111101";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111110111111110";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "0000000011101101";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111010010101";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "0000000011001110";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111010001101";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111001011101";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111001001101";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111111010011110";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111110111000111";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111111001000111";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111000010010";
        wait for Clk_period; 
        Features_din <= "1111111001010110";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111001110100";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111000110101";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111000111111";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111010001111";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "1111111010100100";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111001110001";
        wait for Clk_period; 
        Features_din <= "1111111001011001";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111010011111";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111001111010";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111010001101";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111001111111";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000001001010100";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "0000000011010101";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111011001011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "1111111001010111";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111010000011";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "0000000011000111";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111001000011";
        wait for Clk_period; 
        Features_din <= "1111111010000111";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111010000111";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111001010100";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111000100110";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111000101101";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111010011010";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "0000000011100010";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111110111110101";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111010010000";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "0000001001011010";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111010011011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110100011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000100011101";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "0000000010101101";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111001011010";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111000110110";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111000110100";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000100000111";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "0000000010110011";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "0000000011011110";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111001111011";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111000101001";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111010011111";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111001101110";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111000111011";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111110111011010";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111001111011";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111010011000";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111001011110";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "0000000010111000";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "0000000011110101";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000101001011";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "0000000100000010";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111111010010001";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111001010101";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "0000001001001010";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "0000000011100111";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "1111111001000111";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111101111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010100000";
        wait for Clk_period; 
        Features_din <= "1111111000110100";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000000010111110";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "0000000011101000";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "0000000100101101";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111010011010";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111001100111";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111001110011";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111001101011";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "0000000011100010";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111001101111";
        wait for Clk_period; 
        Features_din <= "1111111001110001";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111000101101";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "0000000011110010";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111001111110";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111010010111";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "0000000011110000";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000000011110111";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111001011101";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111001010000";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111110111111110";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111010011110";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111010101110";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111010101110";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111001101110";
        wait for Clk_period; 
        Features_din <= "1111111001011110";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "1111111001110000";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "0000000100010000";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111010011001";
        wait for Clk_period; 
        Features_din <= "1111111010101000";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111010011111";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111001111101";
        wait for Clk_period; 
        Features_din <= "1111111010001101";
        wait for Clk_period; 
        Features_din <= "1111111001101011";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "0000001100001100";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101110110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010110011";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "0000000010111110";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "1111111000010000";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111010100101";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "0000000011100110";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111000111011";
        wait for Clk_period; 
        Features_din <= "1111111000101101";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "0000000011110101";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111001001111";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111000000001";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111001110100";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111000101110";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111001101000";
        wait for Clk_period; 
        Features_din <= "1111111001011010";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111110111111010";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111001000101";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "0000000101011010";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111010101000";
        wait for Clk_period; 
        Features_din <= "1111111001000011";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111111010001100";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "0000001001000100";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111010100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111001011010";
        wait for Clk_period; 
        Features_din <= "1111111010000000";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "0000000011000110";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "0000000100000001";
        wait for Clk_period; 
        Features_din <= "0000000010110011";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111001111010";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "1111111010000111";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111001101000";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "0000000011100011";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111010001101";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111010001001";
        wait for Clk_period; 
        Features_din <= "1111111000011100";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111000000101";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111010001101";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111001011110";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111000100101";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111010000010";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111010001110";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111001001001";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111000111000";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000011001101";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111001100110";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "1111111010011111";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "0000001010001011";
        wait for Clk_period; 
        Features_din <= "1111111010011011";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "0000000011001100";
        wait for Clk_period; 
        Features_din <= "0000000100001111";
        wait for Clk_period; 
        Features_din <= "1111111010000001";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(5, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101010010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111001011110";
        wait for Clk_period; 
        Features_din <= "1111111010000111";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "0000000100010001";
        wait for Clk_period; 
        Features_din <= "0000000011101100";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111010100000";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "0000000011010111";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "0000000011110110";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111010100000";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111001000010";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "0000000110000110";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "1111111000010111";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111001100000";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000011110110";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111010011011";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111001101101";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111001101100";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111001011001";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111010010101";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111010001101";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111001011000";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111000111110";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111001110011";
        wait for Clk_period; 
        Features_din <= "1111111000111101";
        wait for Clk_period; 
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "0000000011000111";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111010000000";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "0000001100100111";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "1111111001111010";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111100100110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111001110011";
        wait for Clk_period; 
        Features_din <= "1111111001110101";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111000111010";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "0000000011001100";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111010101010";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111001001111";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111001111001";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111010000010";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "0000000010111111";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111000110001";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111010010000";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "0000000011110010";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111010100000";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111010110011";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111110111001010";
        wait for Clk_period; 
        Features_din <= "1111111001101101";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111110111000101";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000001000000111";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111010000010";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101100101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111010110011";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "0000000011110110";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111000001101";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111000111110";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "0000000100100000";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111010000010";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "0000000100011011";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111010011011";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111001101000";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111001001001";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111001000110";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111110111110010";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111001111111";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111000110101";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "1111111010100100";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111000000001";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111000000000";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111010100101";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111001011010";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111000011110";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000011010010";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111000111000";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111000110001";
        wait for Clk_period; 
        Features_din <= "1111111010011110";
        wait for Clk_period; 
        Features_din <= "1111111010001110";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "0000001001000000";
        wait for Clk_period; 
        Features_din <= "1111111001010011";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000000011010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "0000000011001110";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "0000000011100010";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111001001110";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111010100100";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "0000000100100111";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111001100000";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111000001011";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "0000000010111111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "1111111001101100";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "0000000011001101";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000000101001010";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111000001010";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111010001001";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111001000100";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111010000110";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111001100101";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000100011100";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111001000111";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111010011011";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111010000100";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "0000001001110100";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111010011000";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "0000000011001001";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101011110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111001000110";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "0000000011011110";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111111001111101";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111000001001";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "0000000011001110";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "0000000011110100";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111010001100";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "0000000101111001";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111001011011";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111010011011";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111001011110";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111001011100";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111001001000";
        wait for Clk_period; 
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "1111111000011000";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "0000000010111101";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "0000000100010010";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111001111001";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111010101110";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111010001100";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111000011101";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111001110101";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "1111111010011110";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111010001011";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "0000001001001001";
        wait for Clk_period; 
        Features_din <= "1111111001111001";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(3, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111100111000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111010110011";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "0000000011010010";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111000101010";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111000100100";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111010001101";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111001011000";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111010011001";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111010101000";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "0000000010101100";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111010000100";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111010000110";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111000101010";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "0000000011000111";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111000110011";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111111010011111";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111001110001";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "0000001000000111";
        wait for Clk_period; 
        Features_din <= "1111111000010010";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110111011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111010011010";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "0000000011111011";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111001110011";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "1111111010100100";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "0000000011100010";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "0000000011100001";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "0000000011010001";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "0000000011110001";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111000101111";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "0000000011011000";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111001100111";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111000011011";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "0000000101000010";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111000010101";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111010101000";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111001011011";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111001011101";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "0000000011101101";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111001010100";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111010001100";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "0000000100100011";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "0000000011000100";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "0000000111001011";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111001110000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110110100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111001011000";
        wait for Clk_period; 
        Features_din <= "1111111001000011";
        wait for Clk_period; 
        Features_din <= "1111111010001111";
        wait for Clk_period; 
        Features_din <= "0000000011101110";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111110111110111";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111001100001";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111010100101";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111010010011";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "0000000110010011";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111110111001111";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111010100100";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111001111100";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111010000001";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000010101100";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "1111111001010001";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "0000000010111100";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111001010100";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111010000110";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "0000000101101111";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111010011001";
        wait for Clk_period; 
        Features_din <= "1111111010001010";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "0000000011010000";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111111010100101";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "1111111001111110";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "0000001100011011";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111100001110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111001011110";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111001001011";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111001101010";
        wait for Clk_period; 
        Features_din <= "1111111010011011";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111010011110";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "0000000011011000";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111001111100";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111000001000";
        wait for Clk_period; 
        Features_din <= "1111111010100000";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111010011001";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111010011000";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111010011011";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111000110000";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111001111011";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111001100001";
        wait for Clk_period; 
        Features_din <= "1111111001001001";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "0000000101111100";
        wait for Clk_period; 
        Features_din <= "1111110111011101";
        wait for Clk_period; 
        Features_din <= "1111111001110100";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101000100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111001011000";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "0000000100000101";
        wait for Clk_period; 
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111001101111";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111010010101";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111001111111";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "1111111001101101";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111010100101";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111001001000";
        wait for Clk_period; 
        Features_din <= "1111111000110000";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111000000010";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111010011001";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111001000101";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111010011110";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "0000000011100100";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111001101110";
        wait for Clk_period; 
        Features_din <= "1111111001110111";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "0000000011100000";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000011100111";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "0000000011010011";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111000110100";
        wait for Clk_period; 
        Features_din <= "1111110111111101";
        wait for Clk_period; 
        Features_din <= "1111111001101000";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000001001110010";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000000011111110";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111001111011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101000000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111001001001";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "1111111001110010";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111111010001010";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "0000000100101100";
        wait for Clk_period; 
        Features_din <= "1111111010101000";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000000011010010";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111001001101";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111010011110";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111010000111";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "0000000100010011";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111110111111001";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "0000000011010010";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111001111000";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "0000000011100010";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111010010111";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111000110101";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111010001100";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "0000000011001111";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "0000000011000111";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "1111111001010111";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111110110101100";
        wait for Clk_period; 
        Features_din <= "1111111010100101";
        wait for Clk_period; 
        Features_din <= "1111111001011100";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111001101110";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "0000000111010011";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111010000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111111001010100";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "0000000100011010";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111000110011";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111010001111";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111000111000";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "0000000100001110";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111001100100";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111110111110110";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111010010111";
        wait for Clk_period; 
        Features_din <= "1111111001111101";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "0000000100010000";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "0000000010101101";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111001101001";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111110111101110";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111010011111";
        wait for Clk_period; 
        Features_din <= "1111111010011111";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "0000001000000101";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111000011001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110011010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111001010111";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "0000000011111000";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111001110001";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111001100001";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "0000000100100001";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "0000000011010010";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111001111111";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "0000000100110010";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111001011010";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111001110100";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111010010000";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111001111111";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111001010010";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111001111010";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111001000100";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111010010101";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111110110011010";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111001111111";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111010011110";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111000011111";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000000100001000";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "1111111001110111";
        wait for Clk_period; 
        Features_din <= "1111111001011100";
        wait for Clk_period; 
        Features_din <= "1111111010000000";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "0000001011111010";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "0000000011100101";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111100110000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111010001001";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111111000101100";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111010110011";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "0000000100011010";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111010101010";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111001110001";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "0000000100011101";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "0000000010111000";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111001010011";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111001110011";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111010001111";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111010000010";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111001001111";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "0000000010111101";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "1111111001110101";
        wait for Clk_period; 
        Features_din <= "1111111010011111";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "0000000110101001";
        wait for Clk_period; 
        Features_din <= "1111111010001011";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "1111111001110011";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110010111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010010111";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000011011011";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "0000000100010010";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "1111111010010101";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111001110010";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111000111111";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111001110011";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "0000000011011110";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111000100100";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "0000000011110110";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111110111011101";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "0000000011001101";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111001110111";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111001011100";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "0000000100110101";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111001110111";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111111000101000";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111000000101";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111001011101";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111001110000";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111001100110";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111010000111";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111001110101";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "0000000011000100";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111001111000";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000000100010001";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111010001101";
        wait for Clk_period; 
        Features_din <= "1111111001000010";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "1111111010000100";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "0000001001000010";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111111010011010";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111100001110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111001001010";
        wait for Clk_period; 
        Features_din <= "1111111010100100";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "0000000010111100";
        wait for Clk_period; 
        Features_din <= "0000000011111001";
        wait for Clk_period; 
        Features_din <= "1111111010001001";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111001010100";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111000101001";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111001111011";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111010010101";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111001000101";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111000101001";
        wait for Clk_period; 
        Features_din <= "1111111000111000";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111110110001100";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "1111111001010101";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111001001011";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "0000000011001110";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111010100000";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111000110101";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111010100101";
        wait for Clk_period; 
        Features_din <= "1111111001111101";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111001000010";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000011100111";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000011100000";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111001000010";
        wait for Clk_period; 
        Features_din <= "1111110111111000";
        wait for Clk_period; 
        Features_din <= "1111111000110110";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111010010111";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "0000001010110111";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "0000000011000101";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111100010111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111010000000";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111000001110";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111001110111";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111001011110";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111010001010";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111010011001";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000010101100";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111000010000";
        wait for Clk_period; 
        Features_din <= "1111111001000000";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "0000000011001010";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "0000000100110000";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111001111111";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000000011010010";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111001101010";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111010100100";
        wait for Clk_period; 
        Features_din <= "1111111000101011";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "1111111000000011";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "0000000010110011";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101010100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111000101101";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "0000000100010000";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111001110001";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111000111011";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111010000110";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111001010101";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "0000000011010001";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111010011001";
        wait for Clk_period; 
        Features_din <= "1111111010010000";
        wait for Clk_period; 
        Features_din <= "1111111001001111";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "0000000100010011";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111001111010";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111001011111";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111010000111";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111001111100";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "0000000011110111";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111110111010110";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111010101000";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111010011010";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111000000111";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111001101001";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111010011110";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111010001110";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000100000100";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "0000000011100011";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111001101010";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111010011011";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111001111101";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "0000000111001101";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "0000000011100001";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101110000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "1111111001000111";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "0000000010110011";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111000000011";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111001001011";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "0000000011001011";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111001111110";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111001110011";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111010001011";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "1111111001111011";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111000111111";
        wait for Clk_period; 
        Features_din <= "1111111010011111";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111001011110";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111110111011110";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "0000000011011100";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111010001001";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111001011010";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111110111111001";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "1111111010000001";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000001010110100";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "0000000010111000";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101101001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111111000011110";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "0000000011010110";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "0000000011101111";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111001011101";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111001011001";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "0000000011101001";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "1111111010000011";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111010011001";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111010000100";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111001011100";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000011111110";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111010011010";
        wait for Clk_period; 
        Features_din <= "1111111010011010";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111110111110111";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "0000000111010011";
        wait for Clk_period; 
        Features_din <= "1111110110010110";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101010111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "0000000011000110";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "0000000101001100";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111010010001";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111010001100";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111010001100";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "0000000100001010";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111001101001";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111000110010";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111001100110";
        wait for Clk_period; 
        Features_din <= "1111111010100100";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111001100100";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111000111101";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111010100000";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111110111010011";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "0000000011010010";
        wait for Clk_period; 
        Features_din <= "0000000011100000";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111001110111";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111001110100";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111010101110";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111010101010";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000001000110011";
        wait for Clk_period; 
        Features_din <= "1111111001011101";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(5, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110010110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111001001010";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111000010111";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "0000000011110001";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "0000000011111101";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111001100110";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111010011110";
        wait for Clk_period; 
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "0000000100000001";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111001010010";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111000000100";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000000010110011";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "1111111010001100";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111000101011";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111001101011";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111001010000";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111000001101";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111010001010";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111010011010";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111000100101";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111110111011110";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111010110011";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "1111111010010001";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111010001001";
        wait for Clk_period; 
        Features_din <= "1111111001011000";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111001110010";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "0000001010011001";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111010101110";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000000100011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111001111100";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "0000000100010000";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111010001011";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "0000000100010110";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "0000000100010100";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111010101010";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "0000000101001000";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111110111001111";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "0000000011010000";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "0000000010101101";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111001110111";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111111000001001";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "0000000101011001";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111010010111";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111001101000";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111010000001";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000011111111";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111001100110";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111000110000";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "0000001001010011";
        wait for Clk_period; 
        Features_din <= "1111111000000111";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111011111000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111010000111";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111001010101";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "0000000011110110";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111001010010";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "1111111010000100";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111010011110";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "0000000010110010";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111001111000";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111010101010";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "0000000011100000";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111010001111";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111000100001";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "0000000110100011";
        wait for Clk_period; 
        Features_din <= "1111111000010100";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111011001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000011011100";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111001001010";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "0000000011010000";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111010110011";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "0000000100000001";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111010101110";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "0000000011110011";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111010011011";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "0000000011111110";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111001000000";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111001100000";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111010101010";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111000101001";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "0000000101000100";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111010001010";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111001111010";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000001010100100";
        wait for Clk_period; 
        Features_din <= "1111110110101001";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "0000000011101001";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(6, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111100000100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111000101111";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000011010101";
        wait for Clk_period; 
        Features_din <= "1111110111110100";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000011100010";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "0000000010111000";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "1111111001010101";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111010001110";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "0000000010110011";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111001011110";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111010011000";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111010010001";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000011011001";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111111010000110";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111001110111";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "0000000011000100";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111001110001";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "1111111011001110";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111010010101";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111001001000";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "0000001000101001";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111001100100";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110010100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111001110001";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "0000000011101101";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "1111111001101001";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111000101000";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111110111110111";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "0000000011111111";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111000110111";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000011100110";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "0000000011000001";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111001001110";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "0000000101110101";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111000001000";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111000100101";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111001100000";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111010011010";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111010001100";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111110111111111";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111001111111";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111001010011";
        wait for Clk_period; 
        Features_din <= "1111111010001010";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111001011011";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111001101001";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111010001011";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111001101111";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000000101011110";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "0000000101111001";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111001110000";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111001111110";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "0000001011110011";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101100100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111001110010";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111001110001";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "0000000100111001";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "0000000011000111";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111001111001";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "0000000011011110";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111010000110";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "0000000100100110";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111010010011";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111001000100";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111010010011";
        wait for Clk_period; 
        Features_din <= "1111111001010101";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111110111100101";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "0000000011010010";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111010000110";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "0000001000101000";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101100001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010011000";
        wait for Clk_period; 
        Features_din <= "1111111001010111";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111111010010001";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "0000000101010001";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111001110001";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "0000000010110010";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111010000100";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111010001011";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111001100001";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111000010001";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111000001000";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111010001111";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111001011111";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111001110000";
        wait for Clk_period; 
        Features_din <= "1111111000101010";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "0000001000111011";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111011111011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111000111010";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111001111111";
        wait for Clk_period; 
        Features_din <= "0000000101001111";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111110111111011";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111010001110";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111000111010";
        wait for Clk_period; 
        Features_din <= "1111111001001011";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111001100101";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111010001111";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111010100100";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111010011010";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111010001011";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111111010101000";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111001001010";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111001000011";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111010001011";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111001010001";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "1111111010101000";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111000001011";
        wait for Clk_period; 
        Features_din <= "0000000011101110";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111010000000";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111001110101";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "0000000100111100";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110101000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010001110";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000011001100";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "1111111001011111";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111001011110";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111000110001";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "0000000011100001";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111001111110";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111001111001";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111010010011";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111000011100";
        wait for Clk_period; 
        Features_din <= "1111111001100001";
        wait for Clk_period; 
        Features_din <= "1111111001100011";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111000100001";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "0000000011001000";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111010000000";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000100001111";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111000001000";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111000010001";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "1111110111111111";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111000001010";
        wait for Clk_period; 
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "1111111010101000";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111000011000";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111001110101";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111001100100";
        wait for Clk_period; 
        Features_din <= "1111111000111110";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111001010111";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000101000000";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111010000110";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111001110000";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111001011011";
        wait for Clk_period; 
        Features_din <= "1111111000011100";
        wait for Clk_period; 
        Features_din <= "1111111001001100";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111110111110100";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "0000001000001100";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000011010010";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111001001100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110000111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111001001001";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111001000000";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "0000001000011111";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111000101011";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111010100101";
        wait for Clk_period; 
        Features_din <= "1111111010001011";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111001111001";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111001011001";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111010101010";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111010000000";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111001111101";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111000011001";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111000100001";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111001011100";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111010101110";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "0000000110100101";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "1111111000011100";
        wait for Clk_period; 
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101110010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111001011001";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111001010011";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111010001110";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111000100100";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "0000000011011000";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000101010010";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111010011011";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111001100101";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111010100100";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111111001111101";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111010000110";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "0000000011010001";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111010011001";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111001101001";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111000110100";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111010100000";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111001110001";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111001101000";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "0000000100110101";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111001110101";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111010011110";
        wait for Clk_period; 
        Features_din <= "1111111001010111";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111010010011";
        wait for Clk_period; 
        Features_din <= "0000000010101101";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111001001110";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111010001001";
        wait for Clk_period; 
        Features_din <= "1111111010101010";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111001101010";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "0000001010100110";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "0000000100100010";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(5, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111011000010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111001100001";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "0000000010111101";
        wait for Clk_period; 
        Features_din <= "1111111000110110";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111010001101";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111001011111";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000011001010";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111010001111";
        wait for Clk_period; 
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111111000110111";
        wait for Clk_period; 
        Features_din <= "1111111001101011";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "1111110111000011";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111001111000";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111010001100";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111111001001100";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "1111111001101010";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111000101100";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "1111111001100110";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111000111010";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111001010001";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111110111110100";
        wait for Clk_period; 
        Features_din <= "1111111001011101";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "0000000011100110";
        wait for Clk_period; 
        Features_din <= "0000000110110111";
        wait for Clk_period; 
        Features_din <= "1111111001110111";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111100110111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111001111101";
        wait for Clk_period; 
        Features_din <= "1111111010000001";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "0000000011111001";
        wait for Clk_period; 
        Features_din <= "0000000011000001";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000011001100";
        wait for Clk_period; 
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111010100010";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111010001100";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111000110001";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111001110000";
        wait for Clk_period; 
        Features_din <= "1111111000000100";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111000001101";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "0000000011000100";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111010111110";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111110111100111";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111110110101001";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111010010111";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "1111111001000001";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111111001001";
        wait for Clk_period; 
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111000011000";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "0000000011010001";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111010000110";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "1111111000110101";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111001110110";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "0000001010101100";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111001111011";
        wait for Clk_period; 
        Features_din <= "0000000011010011";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(6, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110010110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111001111110";
        wait for Clk_period; 
        Features_din <= "1111111000001010";
        wait for Clk_period; 
        Features_din <= "0000000011011110";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111000101011";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111010010111";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "0000000011101011";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111010001110";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111110111111011";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000011101110";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111010011001";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111001110010";
        wait for Clk_period; 
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "0000000100110011";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "0000000011111100";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111001000010";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "0000000011000111";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111001110101";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111000111100";
        wait for Clk_period; 
        Features_din <= "1111111010001001";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "1111111011111100";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111001000000";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111010011011";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000100100111";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "1111111010010000";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "0000000111101110";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111001000110";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111001000010";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "0000001100101011";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110000000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111000110010";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "0000000011000111";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "1111111110100100";
        wait for Clk_period; 
        Features_din <= "1111111010011011";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111001010100";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111111000011";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111001110101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111010100100";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111001101100";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111010110011";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111001100100";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "0000000011000000";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "0000000011011001";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111111010101110";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111111010000001";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111010111000";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111010010000";
        wait for Clk_period; 
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111001000110";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "0000000011110011";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111001011101";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111110010010";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111100011011";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "0000000011010000";
        wait for Clk_period; 
        Features_din <= "0000000011101011";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111010100101";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000000100000010";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111001110011";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "0000001100101001";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111100000110";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111100100011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111000000010";
        wait for Clk_period; 
        Features_din <= "1111111010011111";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "1111111000010011";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111001110101";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111000101111";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "0000000100000100";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111001011101";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111001011111";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "1111111000111110";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111010000011";
        wait for Clk_period; 
        Features_din <= "0000000100111001";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111010001011";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111010000100";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111001011111";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111000110111";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111101000101";
        wait for Clk_period; 
        Features_din <= "1111111110010110";
        wait for Clk_period; 
        Features_din <= "1111111010110101";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111000101111";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111001011111";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111110110000";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111000100100";
        wait for Clk_period; 
        Features_din <= "1111111011111010";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111001110111";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "0000000011000111";
        wait for Clk_period; 
        Features_din <= "0000000011000110";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "1111111001001111";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "1111111001110010";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111111100001";
        wait for Clk_period; 
        Features_din <= "1111111001011110";
        wait for Clk_period; 
        Features_din <= "1111111001001001";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "1111111010001011";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "0000001001100000";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "0000000010111000";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111001111000";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111110010101";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111011111001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111001111100";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000011011101";
        wait for Clk_period; 
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111000001100";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "0000000011100000";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111001111111";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "1111111010011000";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111010100000";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "0000000010111000";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "1111111001001100";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111010000010";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "0000000100100111";
        wait for Clk_period; 
        Features_din <= "1111111110100011";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111101011001";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111110111000110";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "1111111001100110";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "0000000100111001";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111001000100";
        wait for Clk_period; 
        Features_din <= "0000000010111100";
        wait for Clk_period; 
        Features_din <= "1111111001101100";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "1111111011000000";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111010100011";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111101101111";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111100001101";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "0000000011011011";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111111001101101";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "0000000010101100";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111001000111";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111010010101";
        wait for Clk_period; 
        Features_din <= "1111111010001111";
        wait for Clk_period; 
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000010111100";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "1111111001010101";
        wait for Clk_period; 
        Features_din <= "1111111010011001";
        wait for Clk_period; 
        Features_din <= "1111111001011110";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "0000001000001110";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(5, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111101010001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111010010010";
        wait for Clk_period; 
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "0000000100000101";
        wait for Clk_period; 
        Features_din <= "0000000011001011";
        wait for Clk_period; 
        Features_din <= "1111111001110011";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "1111111001001010";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111000001111";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "1111111010011001";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111001101011";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111010001111";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111100000011";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "0000000101101001";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111010001011";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "1111111101011110";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111001111001";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111110000100";
        wait for Clk_period; 
        Features_din <= "1111111101111011";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "1111111101010000";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111110001010";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111100000100";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111001110011";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111010101011";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111000100000";
        wait for Clk_period; 
        Features_din <= "1111111011000101";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "1111111001111000";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111010000000";
        wait for Clk_period; 
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111001001111";
        wait for Clk_period; 
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "1111111101101101";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111101111110";
        wait for Clk_period; 
        Features_din <= "1111111010000010";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111010001110";
        wait for Clk_period; 
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "1111110111001000";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111010000110";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "0000000011001100";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "0000000010111110";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000011001100";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111111110000110";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111010001100";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111001101010";
        wait for Clk_period; 
        Features_din <= "1111111001100110";
        wait for Clk_period; 
        Features_din <= "1111111010100101";
        wait for Clk_period; 
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111110110100";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111101110001";
        wait for Clk_period; 
        Features_din <= "1111111101111010";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111111110100110";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "1111111010110000";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "0000001010110111";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111110001011";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111101110100";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110100000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010010100";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "0000000011010110";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111010010011";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111010000001";
        wait for Clk_period; 
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "1111111001011110";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111001110011";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111101110011";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111001110010";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111111101100011";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111110001101";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "0000000101001011";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "1111111101101011";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111001101001";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111101110101";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111110001111";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111001111100";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111111010010111";
        wait for Clk_period; 
        Features_din <= "1111111010001001";
        wait for Clk_period; 
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "1111111101111001";
        wait for Clk_period; 
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111110011101";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "1111111101100010";
        wait for Clk_period; 
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111111001000111";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111111101001000";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111110011010";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "1111111000010100";
        wait for Clk_period; 
        Features_din <= "1111111100111001";
        wait for Clk_period; 
        Features_din <= "1111111101111101";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111101100100";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "0000000010101101";
        wait for Clk_period; 
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000010111111";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "1111111000100110";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "1111111100011111";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111110011000";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "1111111111001111";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111001110000";
        wait for Clk_period; 
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111101101100";
        wait for Clk_period; 
        Features_din <= "1111111110011011";
        wait for Clk_period; 
        Features_din <= "1111111110010111";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "1111111110000010";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111110100111";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "1111111110001100";
        wait for Clk_period; 
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111010100111";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111101010111";
        wait for Clk_period; 
        Features_din <= "1111111110101000";
        wait for Clk_period; 
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111010100100";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111111110011100";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "1111111011000110";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "1111111101111000";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111010001000";
        wait for Clk_period; 
        Features_din <= "1111111110111010";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "1111111111000010";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111111001110011";
        wait for Clk_period; 
        Features_din <= "1111111110000000";
        wait for Clk_period; 
        Features_din <= "1111111110100101";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000100001001";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111111101101001";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111001101001";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "1111111101101110";
        wait for Clk_period; 
        Features_din <= "1111111010110100";
        wait for Clk_period; 
        Features_din <= "1111111000111110";
        wait for Clk_period; 
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "1111111110111110";
        wait for Clk_period; 
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "1111111001110101";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111110101101";
        wait for Clk_period; 
        Features_din <= "0000001011011101";
        wait for Clk_period; 
        Features_din <= "1111111011011101";
        wait for Clk_period; 
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
            wait;
    end process;
end;
