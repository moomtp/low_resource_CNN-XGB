

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.types.all;

entity image_test is
    generic(TREE_RAM_BITS: positive := 13;
            NUM_CLASSES:   positive := 8;
            NUM_FEATURES:  positive := 35);
end image_test;

architecture behavior of image_test is
    
    component image
        generic(TREE_RAM_BITS: positive;
                NUM_CLASSES:   positive;
                NUM_FEATURES:  positive);
        port(-- Control signals
             Clk:   in std_logic;
             Reset: in std_logic;
             
             -- Inputs for the nodes reception (trees)
             Load_trees: in std_logic;
             Valid_node: in std_logic;
             Addr:       in std_logic_vector(TREE_RAM_BITS - 1  downto 0);
             Trees_din:  in std_logic_vector(31 downto 0);
             
             -- Inputs for the features reception (pixels)
             Load_features: in std_logic;
             Valid_feature: in std_logic;
             Features_din:  in std_logic_vector(15 downto 0);
             Last_feature:  in std_logic;
             
             -- Output signals
             --     Finish:     finish (also 'ready') signal
             --     Dout:       the selected class
             --     Greater:    the value of the selected class prediction
             --     Curr_state: the current state
             Finish:     out std_logic;
             Dout:       out std_logic_vector(log_2(NUM_CLASSES) - 1 downto 0);
             greater:    out std_logic_vector(31 downto 0);
             curr_state: out std_logic_vector(2 downto 0));
    end component;
    
    component counter is
        generic(BITS: natural);
        port(Clk:   in  std_logic;
             Reset: in  std_logic;
             Count: in  std_logic;
             Dout:  out std_logic_vector (BITS - 1 downto 0));
    end component;
    
    -- Inputs
    signal Clk:           std_logic := '0';
    signal Reset:         std_logic := '0';
    signal Load_trees:    std_logic := '0';
    signal Valid_node:    std_logic := '0';
    signal Addr:          std_logic_vector(TREE_RAM_BITS - 1 downto
                                           0) := (others => '0');
    signal Trees_din:     std_logic_vector(31 downto 0) := (others => '0');
    signal Load_features: std_logic := '0';
    signal Valid_feature: std_logic := '0';
    signal Features_din:  std_logic_vector(15 downto 0) := (others => '0');
    signal last_feature:  std_logic := '0';
    
    -- Outputs
    signal Finish:     std_logic;
    signal Dout:       std_logic_vector(log_2(NUM_CLASSES) - 1 downto 0);
    signal greater:    std_logic_vector(31 downto 0);
    signal curr_state: std_logic_vector(2 downto 0);
    
    -- Clock period definition
    constant Clk_period : time := 10 ns;
    
    -- Counter signals
    signal pc_count, hc_count: std_logic := '0';
    signal pixels, hits: std_logic_vector(15 downto 0) := (others => '0');
    
    -- Label signal
    signal class_label: std_logic_vector(log_2(NUM_CLASSES) - 1 downto 0);

begin
    
    -- Instantiate the Unit Under Test (UUT)
    uut: image
        generic map(TREE_RAM_BITS => TREE_RAM_BITS,
                    NUM_CLASSES   => NUM_CLASSES,
                    NUM_FEATURES  => NUM_FEATURES)
        port map(Clk           => Clk,
                 Reset         => Reset,
                 Load_trees    => Load_trees,
                 Valid_node    => Valid_node,
                 Addr          => Addr,
                 Trees_din     => Trees_din,
                 Load_features => Load_features,
                 Valid_feature => Valid_feature,
                 Features_din  => Features_din,
                 Last_feature  => Last_feature,
                 Finish        => Finish,
                 Dout          => Dout,
                 greater       => greater,
                 curr_state    => curr_state);
    
    -- To count the pixels
    pixel_counter: counter
        generic map(BITS => 16)
        port map(Clk   => Clk, 
                 Reset => Reset,
                 Count => pc_count,
                 Dout  => pixels);
    
    -- To count the hits
    hit_counter: counter
        generic map(BITS => 16)
        port map(Clk   => Clk, 
                 Reset => Reset,
                 Count => hc_count,
                 Dout  => hits);
    
    -- Clock process definition
    Clk_process: process
    begin
        Clk <= '0';
        wait for Clk_period/2;
        Clk <= '1';
        wait for Clk_period/2;
    end process;
    
    -- Stimulus process
    stim_proc: process
    begin
        
        Reset <= '1';
        
        -- hold reset state for 100 ns.
        wait for 100 ns;
        
        Reset <= '0';
        
        wait for Clk_period*10;
        


        
        -- LOAD TREES
        -----------------------------------------------------------------------
        
        -- Load and valid trees flags
        Load_trees <= '1';
        Valid_node <= '1';

        -- Class  0
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"06082678";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"0605c338";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"06038618";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"06005808";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"14005904";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"ff540195";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"00000195";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"08005608";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"00fe7704";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"ff550195";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"ff970195";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"08005804";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"015c0195";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"ff7c0195";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"00ff0810";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"09003708";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"00fd3704";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"ffa70195";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"01660195";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"1f028204";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"ff8a0195";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"00570195";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"09003c08";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"0e001804";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"00df0195";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"ff980195";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"07025c04";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"00230195";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"016e0195";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"04068420";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"03043710";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"0606c708";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"00fe8804";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"014f0195";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"00640195";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"0000da04";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"01f00195";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"00090195";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"15f7ad08";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"05005104";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"01290195";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"ff960195";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"07fe6404";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"ff6a0195";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"00370195";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"01fedd10";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"06077b08";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"18006604";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"ffec0195";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"00ce0195";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"1afe3c04";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"ff750195";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"00ca0195";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"02fb0e08";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"0e002904";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"030e0195";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"00ab0195";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"00fdf404";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"ff900195";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"00370195";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"060a7e2c";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"03067c20";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"04057010";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"04fb9608";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"01fd3304";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"00370195";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"ffa40195";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"0e002304";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"021e0195";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"03490195";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"03feef08";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"0406d404";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"02610195";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"017e0195";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"00fdf604";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"00ca0195";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"ff8c0195";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"0c000704";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"015c0195";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"0307f804";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"00370195";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"ff630195";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"0309a418";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"060b2c0c";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"0305fb08";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"01ffcd04";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"03a40195";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"01290195";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"00c20195";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"05098508";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"0f00a104";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"04680195";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"025f0195";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"00df0195";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"00fd6508";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"0b00ab04";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"00000195";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"02470195";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"00fe7e04";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"ff7e0195";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"00c20195";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"0606d168";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"06040e2c";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"06005810";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"1400590c";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"14003008";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"01fddd04";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"00310321";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"ff620321";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"ff570321";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"000a0321";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"0e002f0c";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"17023108";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"1b027c04";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"003e0321";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"ffa20321";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"ff590321";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"1300b408";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"18006404";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"00900321";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"ff880321";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"00fe6704";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"ffc50321";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"01680321";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"0605c320";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"07025c10";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"01fcf908";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"1000d804";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"ffcf0321";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"018a0321";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"09003704";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"006b0321";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"ff990321";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"1b026608";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"13009e04";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"005b0321";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"ff690321";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"0406e104";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"014d0321";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"fff30321";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"05feaf10";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"02fcec08";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"0b00ed04";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"005d0321";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"01300321";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"0402d004";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"000a0321";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"01d60321";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"19001808";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"0500fe04";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"ff610321";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"004c0321";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"01140321";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"06097734";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"03043720";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"18009410";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"04078108";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"1702cb04";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"00a10321";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"01210321";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"0f008904";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"ffed0321";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"020a0321";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"04068408";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"11003a04";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"021e0321";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"00870321";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"0f005a04";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"ff910321";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"01a90321";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"0c002408";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"05005104";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"018b0321";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"00270321";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"03067c08";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"11000b04";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"ff730321";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"00a50321";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"ff690321";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"030b271c";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"060d3210";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"03067c08";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"04050004";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"01930321";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"014e0321";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"1300a704";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"01340321";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"ffa70321";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"1dfe5e08";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"00fd8a04";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"01070321";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"00050321";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"01c10321";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"02ff5e08";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"17027304";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"00380321";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"ff6c0321";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"0500a704";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"02100321";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"fff00321";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"0605c354";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"06038620";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"06ffb808";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"14005904";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"ff5d047d";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"0022047d";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"19002110";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"02f99f08";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"00ffd204";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"ff6c047d";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"00d4047d";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"06023604";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"ff5d047d";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"ffa2047d";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"0a000b04";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"0152047d";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"ff85047d";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"00ff1d1c";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"0900370c";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"0f008408";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"00fd3704";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"ffd0047d";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"015f047d";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"ff7c047d";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"08005408";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"1af9c104";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"0095047d";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"ff96047d";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"0d008d04";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"0168047d";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"ff84047d";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"05fc1408";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"19000404";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"ff68047d";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"00c7047d";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"05fce508";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"09003604";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"ff93047d";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"0142047d";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"0d006004";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"016e047d";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"ffc1047d";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"0608da2c";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"0406fe18";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"0307f810";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"10034f08";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"05fc2c04";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"0001047d";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"00ba047d";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"02fa2804";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"00d2047d";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"ff7a047d";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"1e024a04";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"0040047d";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"ff72047d";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"01fd4604";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"ff61047d";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"1afcfb08";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"1703e204";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"0044047d";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"0143047d";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"17040004";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"ff5d047d";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"0071047d";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"060c171c";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"03067c10";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"01fc6c08";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"0b00d604";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"00f1047d";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"0049047d";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"0a03b804";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"0107047d";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"0044047d";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"060bac08";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"060abb04";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"ffe0047d";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"0118047d";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"ff62047d";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"030ebc10";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"10000208";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"14003d04";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"ffa0047d";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"0104047d";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"050a7004";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"0132047d";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"001f047d";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"ffa0047d";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"0605334c";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"06038620";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"06ffb808";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"14005904";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"ff6005d9";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"002205d9";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"19002110";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"15f7c808";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"1afcd604";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"002505d9";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"ff6505d9";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"08003c04";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"fff205d9";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"ff5f05d9";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"0a000b04";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"010905d9";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"ff8b05d9";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"02fa3610";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"00ff1204";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"ff6305d9";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"1300a408";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"11000504";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"ffa305d9";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"014205d9";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"ff8405d9";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"0403d20c";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"0603a104";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"008f05d9";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"03071b04";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"ff6305d9";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"003005d9";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"0405d808";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"01fe2b04";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"012d05d9";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"ffe505d9";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"0f007604";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"ff6805d9";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"003d05d9";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"06097738";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"06072d1c";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"0f00870c";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"0f008708";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"1b025404";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"fff805d9";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"006805d9";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"019705d9";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"01fee308";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"16040004";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"ff8405d9";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"00b405d9";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"00fe2704";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"ff8f05d9";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"014d05d9";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"18009410";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"0c02d808";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"03018604";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"009405d9";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"001805d9";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"0f007004";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"00af05d9";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"ff9405d9";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"08005b08";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"03fad104";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"003305d9";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"012b05d9";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"fffc05d9";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"060c1718";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"0306ca0c";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"1af87f04";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"ffb405d9";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"00fdab04";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"00a805d9";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"00d305d9";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"060bac08";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"060aff04";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"ffae05d9";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"00d705d9";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"ff7105d9";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"030ebc10";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"060d6808";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"05063404";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"00e105d9";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"ffc905d9";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"1ffd1c04";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"006605d9";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"010005d9";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"ffa605d9";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"06053360";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"0603862c";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"06ffb810";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"1400590c";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"14002e08";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"17030304";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"003c0775";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"ff780775";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"ff600775";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"00240775";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"19002110";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"02f99f08";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"00ffd204";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"ff770775";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"00d30775";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"06023604";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"ff630775";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"ffb80775";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"0a000b08";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"01fed904";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"01240775";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"00260775";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"ff910775";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"14003b14";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"1400320c";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"06044104";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"ff8a0775";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"04055c04";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"010b0775";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"000a0775";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"01ffbf04";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"ff600775";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"002e0775";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"1300a910";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"03003908";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"00ff2a04";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"ff760775";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"002f0775";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"0b00ec04";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"011d0775";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"ffaa0775";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"12004808";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"05fd0104";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"01860775";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"00100775";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"11004404";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"ffa60775";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"01280775";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"0609e53c";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"01fd091c";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"17023f0c";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"1002e608";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"05ff1c04";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"011c0775";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"fff60775";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"ff820775";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"14004508";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"10000a04";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"ff340775";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"000f0775";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"0a007404";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"00be0775";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"ffb60775";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"10007610";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"1603fd08";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"12003804";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"ffe50775";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"00e40775";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"00fcc204";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"ffdf0775";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"007e0775";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"1603ea08";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"07fed204";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"00210775";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"008a0775";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"14003e04";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"ff9c0775";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"00480775";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"060d3220";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"04fc0c10";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"04fae408";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"ffd80775";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"00b10775";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"19000204";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"ff920775";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"00810775";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"11022308";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"0e005c04";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"00af0775";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"ffbe0775";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"14004804";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"006f0775";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"ff230775";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"01fae008";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"11004704";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"00a10775";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"ffa10775";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"1af87f04";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"00220775";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"04f9fd04";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"009f0775";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"00dd0775";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"06040e34";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"06005810";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"1400590c";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"14003008";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"01fddd04";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"006208c9";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"ff7708c9";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"ff6208c9";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"001d08c9";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"0e002f08";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"05fb3404";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"001208c9";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"ff6308c9";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"1300ab10";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"03fae008";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"04085f04";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"00df08c9";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"ffa508c9";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"10031c04";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"ff7508c9";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"005308c9";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"0c026608";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"10003d04";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"ff9a08c9";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"011208c9";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"ff8908c9";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"060b2c3c";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"0608831c";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"07fea810";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"13007308";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"0c000704";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"003b08c9";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"015808c9";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"13009d04";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"ff7a08c9";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"001208c9";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"1dfd8904";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"ff6108c9";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"05fe1f04";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"005108c9";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"000f08c9";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"01fd0910";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"0b00dc08";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"09004a04";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"008008c9";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"ffa408c9";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"18005704";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"ff4308c9";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"002708c9";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"0305fb08";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"00fd9b04";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"005508c9";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"008c08c9";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"1d024c04";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"00d808c9";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"ff7908c9";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"060d6820";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"0b004b10";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"1602fc08";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"0e002b04";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"00bf08c9";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"ffcc08c9";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"0a00be04";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"002508c9";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"ff2408c9";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"07fc1008";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"10000904";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"ffc708c9";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"007a08c9";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"0b011f04";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"00a908c9";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"ffb008c9";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"04f9fd10";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"060e7708";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"02ff8504";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"ff4b08c9";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"00b908c9";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"030aad04";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"00db08c9";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"ffe008c9";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"0505c808";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"0a000004";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"007508c9";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"00ce08c9";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"000608c9";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"06040e34";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"06ffb810";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"1400590c";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"14002e08";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"0c01c504";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"ff820a1d";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"00430a1d";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"ff640a1d";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"002c0a1d";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"0e002f0c";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"06ffea04";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"002d0a1d";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"17023104";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"00170a1d";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"ff660a1d";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"1300ab0c";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"08004308";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"1703ef04";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"ffa80a1d";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"00ba0a1d";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"ff6c0a1d";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"0c026608";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"02f97104";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"ff960a1d";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"00cc0a1d";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"ff8e0a1d";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"060b2c3c";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"06088320";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"18008e10";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"08004408";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"13009a04";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"ffeb0a1d";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"004d0a1d";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"1d027404";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"ffe70a1d";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"00330a1d";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"11000108";
		wait for Clk_period;
		Addr <=  "0001001010111";
		Trees_din <= x"15f76a04";
		wait for Clk_period;
		Addr <=  "0001001011000";
		Trees_din <= x"00630a1d";
		wait for Clk_period;
		Addr <=  "0001001011001";
		Trees_din <= x"ff640a1d";
		wait for Clk_period;
		Addr <=  "0001001011010";
		Trees_din <= x"10005404";
		wait for Clk_period;
		Addr <=  "0001001011011";
		Trees_din <= x"01600a1d";
		wait for Clk_period;
		Addr <=  "0001001011100";
		Trees_din <= x"00090a1d";
		wait for Clk_period;
		Addr <=  "0001001011101";
		Trees_din <= x"01fd960c";
		wait for Clk_period;
		Addr <=  "0001001011110";
		Trees_din <= x"0a03c708";
		wait for Clk_period;
		Addr <=  "0001001011111";
		Trees_din <= x"08004a04";
		wait for Clk_period;
		Addr <=  "0001001100000";
		Trees_din <= x"002d0a1d";
		wait for Clk_period;
		Addr <=  "0001001100001";
		Trees_din <= x"00820a1d";
		wait for Clk_period;
		Addr <=  "0001001100010";
		Trees_din <= x"ff250a1d";
		wait for Clk_period;
		Addr <=  "0001001100011";
		Trees_din <= x"0d007208";
		wait for Clk_period;
		Addr <=  "0001001100100";
		Trees_din <= x"11025004";
		wait for Clk_period;
		Addr <=  "0001001100101";
		Trees_din <= x"00910a1d";
		wait for Clk_period;
		Addr <=  "0001001100110";
		Trees_din <= x"ff6a0a1d";
		wait for Clk_period;
		Addr <=  "0001001100111";
		Trees_din <= x"0406fe04";
		wait for Clk_period;
		Addr <=  "0001001101000";
		Trees_din <= x"003a0a1d";
		wait for Clk_period;
		Addr <=  "0001001101001";
		Trees_din <= x"00f70a1d";
		wait for Clk_period;
		Addr <=  "0001001101010";
		Trees_din <= x"060d681c";
		wait for Clk_period;
		Addr <=  "0001001101011";
		Trees_din <= x"07fc1010";
		wait for Clk_period;
		Addr <=  "0001001101100";
		Trees_din <= x"060ce508";
		wait for Clk_period;
		Addr <=  "0001001101101";
		Trees_din <= x"05fe9704";
		wait for Clk_period;
		Addr <=  "0001001101110";
		Trees_din <= x"00d20a1d";
		wait for Clk_period;
		Addr <=  "0001001101111";
		Trees_din <= x"00300a1d";
		wait for Clk_period;
		Addr <=  "0001001110000";
		Trees_din <= x"0e002a04";
		wait for Clk_period;
		Addr <=  "0001001110001";
		Trees_din <= x"ff440a1d";
		wait for Clk_period;
		Addr <=  "0001001110010";
		Trees_din <= x"00690a1d";
		wait for Clk_period;
		Addr <=  "0001001110011";
		Trees_din <= x"0b012708";
		wait for Clk_period;
		Addr <=  "0001001110100";
		Trees_din <= x"08004104";
		wait for Clk_period;
		Addr <=  "0001001110101";
		Trees_din <= x"006a0a1d";
		wait for Clk_period;
		Addr <=  "0001001110110";
		Trees_din <= x"00a10a1d";
		wait for Clk_period;
		Addr <=  "0001001110111";
		Trees_din <= x"ff860a1d";
		wait for Clk_period;
		Addr <=  "0001001111000";
		Trees_din <= x"0305bc10";
		wait for Clk_period;
		Addr <=  "0001001111001";
		Trees_din <= x"0f005708";
		wait for Clk_period;
		Addr <=  "0001001111010";
		Trees_din <= x"10000d04";
		wait for Clk_period;
		Addr <=  "0001001111011";
		Trees_din <= x"00780a1d";
		wait for Clk_period;
		Addr <=  "0001001111100";
		Trees_din <= x"ffd60a1d";
		wait for Clk_period;
		Addr <=  "0001001111101";
		Trees_din <= x"1dfe5e04";
		wait for Clk_period;
		Addr <=  "0001001111110";
		Trees_din <= x"00240a1d";
		wait for Clk_period;
		Addr <=  "0001001111111";
		Trees_din <= x"00be0a1d";
		wait for Clk_period;
		Addr <=  "0001010000000";
		Trees_din <= x"20040008";
		wait for Clk_period;
		Addr <=  "0001010000001";
		Trees_din <= x"08004204";
		wait for Clk_period;
		Addr <=  "0001010000010";
		Trees_din <= x"001d0a1d";
		wait for Clk_period;
		Addr <=  "0001010000011";
		Trees_din <= x"ff3b0a1d";
		wait for Clk_period;
		Addr <=  "0001010000100";
		Trees_din <= x"12003404";
		wait for Clk_period;
		Addr <=  "0001010000101";
		Trees_din <= x"ffaf0a1d";
		wait for Clk_period;
		Addr <=  "0001010000110";
		Trees_din <= x"00b50a1d";
		wait for Clk_period;
		Addr <=  "0001010000111";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0001010001000";
		Trees_din <= x"06040e38";
		wait for Clk_period;
		Addr <=  "0001010001001";
		Trees_din <= x"06ffb810";
		wait for Clk_period;
		Addr <=  "0001010001010";
		Trees_din <= x"1400590c";
		wait for Clk_period;
		Addr <=  "0001010001011";
		Trees_din <= x"14002e08";
		wait for Clk_period;
		Addr <=  "0001010001100";
		Trees_din <= x"0c01c504";
		wait for Clk_period;
		Addr <=  "0001010001101";
		Trees_din <= x"ff880b65";
		wait for Clk_period;
		Addr <=  "0001010001110";
		Trees_din <= x"003d0b65";
		wait for Clk_period;
		Addr <=  "0001010001111";
		Trees_din <= x"ff660b65";
		wait for Clk_period;
		Addr <=  "0001010010000";
		Trees_din <= x"002d0b65";
		wait for Clk_period;
		Addr <=  "0001010010001";
		Trees_din <= x"0e002f0c";
		wait for Clk_period;
		Addr <=  "0001010010010";
		Trees_din <= x"06ffea04";
		wait for Clk_period;
		Addr <=  "0001010010011";
		Trees_din <= x"00310b65";
		wait for Clk_period;
		Addr <=  "0001010010100";
		Trees_din <= x"05fb3404";
		wait for Clk_period;
		Addr <=  "0001010010101";
		Trees_din <= x"00170b65";
		wait for Clk_period;
		Addr <=  "0001010010110";
		Trees_din <= x"ff680b65";
		wait for Clk_period;
		Addr <=  "0001010010111";
		Trees_din <= x"1300ab10";
		wait for Clk_period;
		Addr <=  "0001010011000";
		Trees_din <= x"03fae008";
		wait for Clk_period;
		Addr <=  "0001010011001";
		Trees_din <= x"15f78504";
		wait for Clk_period;
		Addr <=  "0001010011010";
		Trees_din <= x"00df0b65";
		wait for Clk_period;
		Addr <=  "0001010011011";
		Trees_din <= x"ffa90b65";
		wait for Clk_period;
		Addr <=  "0001010011100";
		Trees_din <= x"10031c04";
		wait for Clk_period;
		Addr <=  "0001010011101";
		Trees_din <= x"ff7c0b65";
		wait for Clk_period;
		Addr <=  "0001010011110";
		Trees_din <= x"00500b65";
		wait for Clk_period;
		Addr <=  "0001010011111";
		Trees_din <= x"0c026608";
		wait for Clk_period;
		Addr <=  "0001010100000";
		Trees_din <= x"10003d04";
		wait for Clk_period;
		Addr <=  "0001010100001";
		Trees_din <= x"ff980b65";
		wait for Clk_period;
		Addr <=  "0001010100010";
		Trees_din <= x"00ad0b65";
		wait for Clk_period;
		Addr <=  "0001010100011";
		Trees_din <= x"ff940b65";
		wait for Clk_period;
		Addr <=  "0001010100100";
		Trees_din <= x"060b2c30";
		wait for Clk_period;
		Addr <=  "0001010100101";
		Trees_din <= x"06088318";
		wait for Clk_period;
		Addr <=  "0001010100110";
		Trees_din <= x"0b004b08";
		wait for Clk_period;
		Addr <=  "0001010100111";
		Trees_din <= x"1bfaa804";
		wait for Clk_period;
		Addr <=  "0001010101000";
		Trees_din <= x"001a0b65";
		wait for Clk_period;
		Addr <=  "0001010101001";
		Trees_din <= x"ff600b65";
		wait for Clk_period;
		Addr <=  "0001010101010";
		Trees_din <= x"10007608";
		wait for Clk_period;
		Addr <=  "0001010101011";
		Trees_din <= x"14004a04";
		wait for Clk_period;
		Addr <=  "0001010101100";
		Trees_din <= x"00260b65";
		wait for Clk_period;
		Addr <=  "0001010101101";
		Trees_din <= x"00970b65";
		wait for Clk_period;
		Addr <=  "0001010101110";
		Trees_din <= x"1000d004";
		wait for Clk_period;
		Addr <=  "0001010101111";
		Trees_din <= x"ffba0b65";
		wait for Clk_period;
		Addr <=  "0001010110000";
		Trees_din <= x"002b0b65";
		wait for Clk_period;
		Addr <=  "0001010110001";
		Trees_din <= x"0d00ae10";
		wait for Clk_period;
		Addr <=  "0001010110010";
		Trees_din <= x"03fa7508";
		wait for Clk_period;
		Addr <=  "0001010110011";
		Trees_din <= x"1001d904";
		wait for Clk_period;
		Addr <=  "0001010110100";
		Trees_din <= x"00d20b65";
		wait for Clk_period;
		Addr <=  "0001010110101";
		Trees_din <= x"ff960b65";
		wait for Clk_period;
		Addr <=  "0001010110110";
		Trees_din <= x"03fb0704";
		wait for Clk_period;
		Addr <=  "0001010110111";
		Trees_din <= x"ffe10b65";
		wait for Clk_period;
		Addr <=  "0001010111000";
		Trees_din <= x"00430b65";
		wait for Clk_period;
		Addr <=  "0001010111001";
		Trees_din <= x"1afa6704";
		wait for Clk_period;
		Addr <=  "0001010111010";
		Trees_din <= x"00070b65";
		wait for Clk_period;
		Addr <=  "0001010111011";
		Trees_din <= x"01000b65";
		wait for Clk_period;
		Addr <=  "0001010111100";
		Trees_din <= x"060d681c";
		wait for Clk_period;
		Addr <=  "0001010111101";
		Trees_din <= x"0b004b0c";
		wait for Clk_period;
		Addr <=  "0001010111110";
		Trees_din <= x"02fa5104";
		wait for Clk_period;
		Addr <=  "0001010111111";
		Trees_din <= x"008c0b65";
		wait for Clk_period;
		Addr <=  "0001011000000";
		Trees_din <= x"0c00dd04";
		wait for Clk_period;
		Addr <=  "0001011000001";
		Trees_din <= x"003a0b65";
		wait for Clk_period;
		Addr <=  "0001011000010";
		Trees_din <= x"ff150b65";
		wait for Clk_period;
		Addr <=  "0001011000011";
		Trees_din <= x"00fe6a08";
		wait for Clk_period;
		Addr <=  "0001011000100";
		Trees_din <= x"17040004";
		wait for Clk_period;
		Addr <=  "0001011000101";
		Trees_din <= x"00680b65";
		wait for Clk_period;
		Addr <=  "0001011000110";
		Trees_din <= x"ffec0b65";
		wait for Clk_period;
		Addr <=  "0001011000111";
		Trees_din <= x"0b005604";
		wait for Clk_period;
		Addr <=  "0001011001000";
		Trees_din <= x"ffba0b65";
		wait for Clk_period;
		Addr <=  "0001011001001";
		Trees_din <= x"00970b65";
		wait for Clk_period;
		Addr <=  "0001011001010";
		Trees_din <= x"0305bc10";
		wait for Clk_period;
		Addr <=  "0001011001011";
		Trees_din <= x"0f005708";
		wait for Clk_period;
		Addr <=  "0001011001100";
		Trees_din <= x"01fe6004";
		wait for Clk_period;
		Addr <=  "0001011001101";
		Trees_din <= x"006e0b65";
		wait for Clk_period;
		Addr <=  "0001011001110";
		Trees_din <= x"ffd10b65";
		wait for Clk_period;
		Addr <=  "0001011001111";
		Trees_din <= x"1dfe5e04";
		wait for Clk_period;
		Addr <=  "0001011010000";
		Trees_din <= x"001c0b65";
		wait for Clk_period;
		Addr <=  "0001011010001";
		Trees_din <= x"00b30b65";
		wait for Clk_period;
		Addr <=  "0001011010010";
		Trees_din <= x"20040008";
		wait for Clk_period;
		Addr <=  "0001011010011";
		Trees_din <= x"01fc7404";
		wait for Clk_period;
		Addr <=  "0001011010100";
		Trees_din <= x"ff430b65";
		wait for Clk_period;
		Addr <=  "0001011010101";
		Trees_din <= x"00100b65";
		wait for Clk_period;
		Addr <=  "0001011010110";
		Trees_din <= x"12003404";
		wait for Clk_period;
		Addr <=  "0001011010111";
		Trees_din <= x"ffb00b65";
		wait for Clk_period;
		Addr <=  "0001011011000";
		Trees_din <= x"00a40b65";
		wait for Clk_period;
		Addr <=  "0001011011001";
		Trees_din <= x"06040e30";
		wait for Clk_period;
		Addr <=  "0001011011010";
		Trees_din <= x"06ffb810";
		wait for Clk_period;
		Addr <=  "0001011011011";
		Trees_din <= x"0e00580c";
		wait for Clk_period;
		Addr <=  "0001011011100";
		Trees_din <= x"0c029604";
		wait for Clk_period;
		Addr <=  "0001011011101";
		Trees_din <= x"ff670cc1";
		wait for Clk_period;
		Addr <=  "0001011011110";
		Trees_din <= x"0d008104";
		wait for Clk_period;
		Addr <=  "0001011011111";
		Trees_din <= x"ff8f0cc1";
		wait for Clk_period;
		Addr <=  "0001011100000";
		Trees_din <= x"00380cc1";
		wait for Clk_period;
		Addr <=  "0001011100001";
		Trees_din <= x"00300cc1";
		wait for Clk_period;
		Addr <=  "0001011100010";
		Trees_din <= x"1e025b04";
		wait for Clk_period;
		Addr <=  "0001011100011";
		Trees_din <= x"ff700cc1";
		wait for Clk_period;
		Addr <=  "0001011100100";
		Trees_din <= x"15f7870c";
		wait for Clk_period;
		Addr <=  "0001011100101";
		Trees_din <= x"0d006f08";
		wait for Clk_period;
		Addr <=  "0001011100110";
		Trees_din <= x"05fcd304";
		wait for Clk_period;
		Addr <=  "0001011100111";
		Trees_din <= x"018c0cc1";
		wait for Clk_period;
		Addr <=  "0001011101000";
		Trees_din <= x"00370cc1";
		wait for Clk_period;
		Addr <=  "0001011101001";
		Trees_din <= x"ffa10cc1";
		wait for Clk_period;
		Addr <=  "0001011101010";
		Trees_din <= x"0a02a208";
		wait for Clk_period;
		Addr <=  "0001011101011";
		Trees_din <= x"15f9f504";
		wait for Clk_period;
		Addr <=  "0001011101100";
		Trees_din <= x"ff910cc1";
		wait for Clk_period;
		Addr <=  "0001011101101";
		Trees_din <= x"003f0cc1";
		wait for Clk_period;
		Addr <=  "0001011101110";
		Trees_din <= x"01fd3304";
		wait for Clk_period;
		Addr <=  "0001011101111";
		Trees_din <= x"00f70cc1";
		wait for Clk_period;
		Addr <=  "0001011110000";
		Trees_din <= x"ff900cc1";
		wait for Clk_period;
		Addr <=  "0001011110001";
		Trees_din <= x"060b2c40";
		wait for Clk_period;
		Addr <=  "0001011110010";
		Trees_din <= x"01fd2220";
		wait for Clk_period;
		Addr <=  "0001011110011";
		Trees_din <= x"17035a10";
		wait for Clk_period;
		Addr <=  "0001011110100";
		Trees_din <= x"1f028408";
		wait for Clk_period;
		Addr <=  "0001011110101";
		Trees_din <= x"0a03c704";
		wait for Clk_period;
		Addr <=  "0001011110110";
		Trees_din <= x"006e0cc1";
		wait for Clk_period;
		Addr <=  "0001011110111";
		Trees_din <= x"ff530cc1";
		wait for Clk_period;
		Addr <=  "0001011111000";
		Trees_din <= x"01fcb804";
		wait for Clk_period;
		Addr <=  "0001011111001";
		Trees_din <= x"ff790cc1";
		wait for Clk_period;
		Addr <=  "0001011111010";
		Trees_din <= x"00450cc1";
		wait for Clk_period;
		Addr <=  "0001011111011";
		Trees_din <= x"14004608";
		wait for Clk_period;
		Addr <=  "0001011111100";
		Trees_din <= x"08004f04";
		wait for Clk_period;
		Addr <=  "0001011111101";
		Trees_din <= x"ffef0cc1";
		wait for Clk_period;
		Addr <=  "0001011111110";
		Trees_din <= x"ff6e0cc1";
		wait for Clk_period;
		Addr <=  "0001011111111";
		Trees_din <= x"1f024004";
		wait for Clk_period;
		Addr <=  "0001100000000";
		Trees_din <= x"00f40cc1";
		wait for Clk_period;
		Addr <=  "0001100000001";
		Trees_din <= x"00250cc1";
		wait for Clk_period;
		Addr <=  "0001100000010";
		Trees_din <= x"1b024b10";
		wait for Clk_period;
		Addr <=  "0001100000011";
		Trees_din <= x"01fdad08";
		wait for Clk_period;
		Addr <=  "0001100000100";
		Trees_din <= x"01fd3004";
		wait for Clk_period;
		Addr <=  "0001100000101";
		Trees_din <= x"00b80cc1";
		wait for Clk_period;
		Addr <=  "0001100000110";
		Trees_din <= x"ff7a0cc1";
		wait for Clk_period;
		Addr <=  "0001100000111";
		Trees_din <= x"1cfea904";
		wait for Clk_period;
		Addr <=  "0001100001000";
		Trees_din <= x"ff3e0cc1";
		wait for Clk_period;
		Addr <=  "0001100001001";
		Trees_din <= x"002e0cc1";
		wait for Clk_period;
		Addr <=  "0001100001010";
		Trees_din <= x"10007608";
		wait for Clk_period;
		Addr <=  "0001100001011";
		Trees_din <= x"00fcd704";
		wait for Clk_period;
		Addr <=  "0001100001100";
		Trees_din <= x"fff80cc1";
		wait for Clk_period;
		Addr <=  "0001100001101";
		Trees_din <= x"00600cc1";
		wait for Clk_period;
		Addr <=  "0001100001110";
		Trees_din <= x"1603ea04";
		wait for Clk_period;
		Addr <=  "0001100001111";
		Trees_din <= x"003a0cc1";
		wait for Clk_period;
		Addr <=  "0001100010000";
		Trees_din <= x"ffe30cc1";
		wait for Clk_period;
		Addr <=  "0001100010001";
		Trees_din <= x"060d6820";
		wait for Clk_period;
		Addr <=  "0001100010010";
		Trees_din <= x"08005610";
		wait for Clk_period;
		Addr <=  "0001100010011";
		Trees_din <= x"08004208";
		wait for Clk_period;
		Addr <=  "0001100010100";
		Trees_din <= x"10000504";
		wait for Clk_period;
		Addr <=  "0001100010101";
		Trees_din <= x"ff670cc1";
		wait for Clk_period;
		Addr <=  "0001100010110";
		Trees_din <= x"00490cc1";
		wait for Clk_period;
		Addr <=  "0001100010111";
		Trees_din <= x"09005004";
		wait for Clk_period;
		Addr <=  "0001100011000";
		Trees_din <= x"00800cc1";
		wait for Clk_period;
		Addr <=  "0001100011001";
		Trees_din <= x"ff870cc1";
		wait for Clk_period;
		Addr <=  "0001100011010";
		Trees_din <= x"1b026808";
		wait for Clk_period;
		Addr <=  "0001100011011";
		Trees_din <= x"0e002704";
		wait for Clk_period;
		Addr <=  "0001100011100";
		Trees_din <= x"ffe80cc1";
		wait for Clk_period;
		Addr <=  "0001100011101";
		Trees_din <= x"00990cc1";
		wait for Clk_period;
		Addr <=  "0001100011110";
		Trees_din <= x"0c01e904";
		wait for Clk_period;
		Addr <=  "0001100011111";
		Trees_din <= x"fee70cc1";
		wait for Clk_period;
		Addr <=  "0001100100000";
		Trees_din <= x"00850cc1";
		wait for Clk_period;
		Addr <=  "0001100100001";
		Trees_din <= x"0305bc10";
		wait for Clk_period;
		Addr <=  "0001100100010";
		Trees_din <= x"0f005708";
		wait for Clk_period;
		Addr <=  "0001100100011";
		Trees_din <= x"0e004004";
		wait for Clk_period;
		Addr <=  "0001100100100";
		Trees_din <= x"ffcc0cc1";
		wait for Clk_period;
		Addr <=  "0001100100101";
		Trees_din <= x"00650cc1";
		wait for Clk_period;
		Addr <=  "0001100100110";
		Trees_din <= x"1dfe5e04";
		wait for Clk_period;
		Addr <=  "0001100100111";
		Trees_din <= x"00140cc1";
		wait for Clk_period;
		Addr <=  "0001100101000";
		Trees_din <= x"00ab0cc1";
		wait for Clk_period;
		Addr <=  "0001100101001";
		Trees_din <= x"20040008";
		wait for Clk_period;
		Addr <=  "0001100101010";
		Trees_din <= x"08004204";
		wait for Clk_period;
		Addr <=  "0001100101011";
		Trees_din <= x"00170cc1";
		wait for Clk_period;
		Addr <=  "0001100101100";
		Trees_din <= x"ff580cc1";
		wait for Clk_period;
		Addr <=  "0001100101101";
		Trees_din <= x"12003404";
		wait for Clk_period;
		Addr <=  "0001100101110";
		Trees_din <= x"ffb30cc1";
		wait for Clk_period;
		Addr <=  "0001100101111";
		Trees_din <= x"00920cc1";
		wait for Clk_period;
		Addr <=  "0001100110000";
		Trees_din <= x"060a7e30";
		wait for Clk_period;
		Addr <=  "0001100110001";
		Trees_din <= x"06013014";
		wait for Clk_period;
		Addr <=  "0001100110010";
		Trees_din <= x"09004d10";
		wait for Clk_period;
		Addr <=  "0001100110011";
		Trees_din <= x"1300ce04";
		wait for Clk_period;
		Addr <=  "0001100110100";
		Trees_din <= x"ff670dbd";
		wait for Clk_period;
		Addr <=  "0001100110101";
		Trees_din <= x"0f008508";
		wait for Clk_period;
		Addr <=  "0001100110110";
		Trees_din <= x"02fc7304";
		wait for Clk_period;
		Addr <=  "0001100110111";
		Trees_din <= x"001f0dbd";
		wait for Clk_period;
		Addr <=  "0001100111000";
		Trees_din <= x"00c90dbd";
		wait for Clk_period;
		Addr <=  "0001100111001";
		Trees_din <= x"ff830dbd";
		wait for Clk_period;
		Addr <=  "0001100111010";
		Trees_din <= x"00410dbd";
		wait for Clk_period;
		Addr <=  "0001100111011";
		Trees_din <= x"1d032e14";
		wait for Clk_period;
		Addr <=  "0001100111100";
		Trees_din <= x"00026210";
		wait for Clk_period;
		Addr <=  "0001100111101";
		Trees_din <= x"00fd9808";
		wait for Clk_period;
		Addr <=  "0001100111110";
		Trees_din <= x"08003b04";
		wait for Clk_period;
		Addr <=  "0001100111111";
		Trees_din <= x"00c70dbd";
		wait for Clk_period;
		Addr <=  "0001101000000";
		Trees_din <= x"fff80dbd";
		wait for Clk_period;
		Addr <=  "0001101000001";
		Trees_din <= x"03fe4504";
		wait for Clk_period;
		Addr <=  "0001101000010";
		Trees_din <= x"00360dbd";
		wait for Clk_period;
		Addr <=  "0001101000011";
		Trees_din <= x"00090dbd";
		wait for Clk_period;
		Addr <=  "0001101000100";
		Trees_din <= x"ff6f0dbd";
		wait for Clk_period;
		Addr <=  "0001101000101";
		Trees_din <= x"0d006b04";
		wait for Clk_period;
		Addr <=  "0001101000110";
		Trees_din <= x"002b0dbd";
		wait for Clk_period;
		Addr <=  "0001101000111";
		Trees_din <= x"ff430dbd";
		wait for Clk_period;
		Addr <=  "0001101001000";
		Trees_din <= x"060d682c";
		wait for Clk_period;
		Addr <=  "0001101001001";
		Trees_din <= x"08003b18";
		wait for Clk_period;
		Addr <=  "0001101001010";
		Trees_din <= x"03fcf908";
		wait for Clk_period;
		Addr <=  "0001101001011";
		Trees_din <= x"08003904";
		wait for Clk_period;
		Addr <=  "0001101001100";
		Trees_din <= x"00200dbd";
		wait for Clk_period;
		Addr <=  "0001101001101";
		Trees_din <= x"fe6d0dbd";
		wait for Clk_period;
		Addr <=  "0001101001110";
		Trees_din <= x"15f70d08";
		wait for Clk_period;
		Addr <=  "0001101001111";
		Trees_din <= x"02fc3104";
		wait for Clk_period;
		Addr <=  "0001101010000";
		Trees_din <= x"fffd0dbd";
		wait for Clk_period;
		Addr <=  "0001101010001";
		Trees_din <= x"ff0a0dbd";
		wait for Clk_period;
		Addr <=  "0001101010010";
		Trees_din <= x"1b028404";
		wait for Clk_period;
		Addr <=  "0001101010011";
		Trees_din <= x"00a80dbd";
		wait for Clk_period;
		Addr <=  "0001101010100";
		Trees_din <= x"ffcc0dbd";
		wait for Clk_period;
		Addr <=  "0001101010101";
		Trees_din <= x"12002a04";
		wait for Clk_period;
		Addr <=  "0001101010110";
		Trees_din <= x"ff5d0dbd";
		wait for Clk_period;
		Addr <=  "0001101010111";
		Trees_din <= x"04066f08";
		wait for Clk_period;
		Addr <=  "0001101011000";
		Trees_din <= x"07fc7b04";
		wait for Clk_period;
		Addr <=  "0001101011001";
		Trees_din <= x"00250dbd";
		wait for Clk_period;
		Addr <=  "0001101011010";
		Trees_din <= x"00620dbd";
		wait for Clk_period;
		Addr <=  "0001101011011";
		Trees_din <= x"08004004";
		wait for Clk_period;
		Addr <=  "0001101011100";
		Trees_din <= x"00b20dbd";
		wait for Clk_period;
		Addr <=  "0001101011101";
		Trees_din <= x"ff760dbd";
		wait for Clk_period;
		Addr <=  "0001101011110";
		Trees_din <= x"0305bc10";
		wait for Clk_period;
		Addr <=  "0001101011111";
		Trees_din <= x"13005e04";
		wait for Clk_period;
		Addr <=  "0001101100000";
		Trees_din <= x"001d0dbd";
		wait for Clk_period;
		Addr <=  "0001101100001";
		Trees_din <= x"1ffd1c04";
		wait for Clk_period;
		Addr <=  "0001101100010";
		Trees_din <= x"00080dbd";
		wait for Clk_period;
		Addr <=  "0001101100011";
		Trees_din <= x"05063404";
		wait for Clk_period;
		Addr <=  "0001101100100";
		Trees_din <= x"00a80dbd";
		wait for Clk_period;
		Addr <=  "0001101100101";
		Trees_din <= x"00450dbd";
		wait for Clk_period;
		Addr <=  "0001101100110";
		Trees_din <= x"20040008";
		wait for Clk_period;
		Addr <=  "0001101100111";
		Trees_din <= x"08004204";
		wait for Clk_period;
		Addr <=  "0001101101000";
		Trees_din <= x"00140dbd";
		wait for Clk_period;
		Addr <=  "0001101101001";
		Trees_din <= x"ff640dbd";
		wait for Clk_period;
		Addr <=  "0001101101010";
		Trees_din <= x"12003404";
		wait for Clk_period;
		Addr <=  "0001101101011";
		Trees_din <= x"ffb50dbd";
		wait for Clk_period;
		Addr <=  "0001101101100";
		Trees_din <= x"0b00e904";
		wait for Clk_period;
		Addr <=  "0001101101101";
		Trees_din <= x"009c0dbd";
		wait for Clk_period;
		Addr <=  "0001101101110";
		Trees_din <= x"ffe70dbd";
		wait for Clk_period;
		Addr <=  "0001101101111";
		Trees_din <= x"060c1750";
		wait for Clk_period;
		Addr <=  "0001101110000";
		Trees_din <= x"06013014";
		wait for Clk_period;
		Addr <=  "0001101110001";
		Trees_din <= x"09004d10";
		wait for Clk_period;
		Addr <=  "0001101110010";
		Trees_din <= x"1300ce04";
		wait for Clk_period;
		Addr <=  "0001101110011";
		Trees_din <= x"ff690ef1";
		wait for Clk_period;
		Addr <=  "0001101110100";
		Trees_din <= x"0f008508";
		wait for Clk_period;
		Addr <=  "0001101110101";
		Trees_din <= x"0f007804";
		wait for Clk_period;
		Addr <=  "0001101110110";
		Trees_din <= x"00c30ef1";
		wait for Clk_period;
		Addr <=  "0001101110111";
		Trees_din <= x"00160ef1";
		wait for Clk_period;
		Addr <=  "0001101111000";
		Trees_din <= x"ff890ef1";
		wait for Clk_period;
		Addr <=  "0001101111001";
		Trees_din <= x"003b0ef1";
		wait for Clk_period;
		Addr <=  "0001101111010";
		Trees_din <= x"06069e1c";
		wait for Clk_period;
		Addr <=  "0001101111011";
		Trees_din <= x"05fd4910";
		wait for Clk_period;
		Addr <=  "0001101111100";
		Trees_din <= x"1b025108";
		wait for Clk_period;
		Addr <=  "0001101111101";
		Trees_din <= x"01fe9504";
		wait for Clk_period;
		Addr <=  "0001101111110";
		Trees_din <= x"ff890ef1";
		wait for Clk_period;
		Addr <=  "0001101111111";
		Trees_din <= x"00910ef1";
		wait for Clk_period;
		Addr <=  "0001110000000";
		Trees_din <= x"03fda804";
		wait for Clk_period;
		Addr <=  "0001110000001";
		Trees_din <= x"004b0ef1";
		wait for Clk_period;
		Addr <=  "0001110000010";
		Trees_din <= x"ffdb0ef1";
		wait for Clk_period;
		Addr <=  "0001110000011";
		Trees_din <= x"0e005308";
		wait for Clk_period;
		Addr <=  "0001110000100";
		Trees_din <= x"0d007d04";
		wait for Clk_period;
		Addr <=  "0001110000101";
		Trees_din <= x"ffa30ef1";
		wait for Clk_period;
		Addr <=  "0001110000110";
		Trees_din <= x"00120ef1";
		wait for Clk_period;
		Addr <=  "0001110000111";
		Trees_din <= x"00e90ef1";
		wait for Clk_period;
		Addr <=  "0001110001000";
		Trees_din <= x"0c000610";
		wait for Clk_period;
		Addr <=  "0001110001001";
		Trees_din <= x"0e005008";
		wait for Clk_period;
		Addr <=  "0001110001010";
		Trees_din <= x"00fe4604";
		wait for Clk_period;
		Addr <=  "0001110001011";
		Trees_din <= x"00c10ef1";
		wait for Clk_period;
		Addr <=  "0001110001100";
		Trees_din <= x"00250ef1";
		wait for Clk_period;
		Addr <=  "0001110001101";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "0001110001110";
		Trees_din <= x"00640ef1";
		wait for Clk_period;
		Addr <=  "0001110001111";
		Trees_din <= x"ff5c0ef1";
		wait for Clk_period;
		Addr <=  "0001110010000";
		Trees_din <= x"15f6f908";
		wait for Clk_period;
		Addr <=  "0001110010001";
		Trees_din <= x"04042504";
		wait for Clk_period;
		Addr <=  "0001110010010";
		Trees_din <= x"00460ef1";
		wait for Clk_period;
		Addr <=  "0001110010011";
		Trees_din <= x"ff7b0ef1";
		wait for Clk_period;
		Addr <=  "0001110010100";
		Trees_din <= x"01fd2504";
		wait for Clk_period;
		Addr <=  "0001110010101";
		Trees_din <= x"000b0ef1";
		wait for Clk_period;
		Addr <=  "0001110010110";
		Trees_din <= x"002c0ef1";
		wait for Clk_period;
		Addr <=  "0001110010111";
		Trees_din <= x"0302c124";
		wait for Clk_period;
		Addr <=  "0001110011000";
		Trees_din <= x"16040014";
		wait for Clk_period;
		Addr <=  "0001110011001";
		Trees_din <= x"04066f10";
		wait for Clk_period;
		Addr <=  "0001110011010";
		Trees_din <= x"11025008";
		wait for Clk_period;
		Addr <=  "0001110011011";
		Trees_din <= x"05fd7a04";
		wait for Clk_period;
		Addr <=  "0001110011100";
		Trees_din <= x"003b0ef1";
		wait for Clk_period;
		Addr <=  "0001110011101";
		Trees_din <= x"009a0ef1";
		wait for Clk_period;
		Addr <=  "0001110011110";
		Trees_din <= x"19000604";
		wait for Clk_period;
		Addr <=  "0001110011111";
		Trees_din <= x"00760ef1";
		wait for Clk_period;
		Addr <=  "0001110100000";
		Trees_din <= x"ff980ef1";
		wait for Clk_period;
		Addr <=  "0001110100001";
		Trees_din <= x"ffb10ef1";
		wait for Clk_period;
		Addr <=  "0001110100010";
		Trees_din <= x"08004304";
		wait for Clk_period;
		Addr <=  "0001110100011";
		Trees_din <= x"ff280ef1";
		wait for Clk_period;
		Addr <=  "0001110100100";
		Trees_din <= x"0f006a04";
		wait for Clk_period;
		Addr <=  "0001110100101";
		Trees_din <= x"008c0ef1";
		wait for Clk_period;
		Addr <=  "0001110100110";
		Trees_din <= x"05fefb04";
		wait for Clk_period;
		Addr <=  "0001110100111";
		Trees_din <= x"00050ef1";
		wait for Clk_period;
		Addr <=  "0001110101000";
		Trees_din <= x"ff5e0ef1";
		wait for Clk_period;
		Addr <=  "0001110101001";
		Trees_din <= x"1afc9320";
		wait for Clk_period;
		Addr <=  "0001110101010";
		Trees_din <= x"060e7710";
		wait for Clk_period;
		Addr <=  "0001110101011";
		Trees_din <= x"1603f808";
		wait for Clk_period;
		Addr <=  "0001110101100";
		Trees_din <= x"09004204";
		wait for Clk_period;
		Addr <=  "0001110101101";
		Trees_din <= x"ff6b0ef1";
		wait for Clk_period;
		Addr <=  "0001110101110";
		Trees_din <= x"001d0ef1";
		wait for Clk_period;
		Addr <=  "0001110101111";
		Trees_din <= x"04fee304";
		wait for Clk_period;
		Addr <=  "0001110110000";
		Trees_din <= x"00940ef1";
		wait for Clk_period;
		Addr <=  "0001110110001";
		Trees_din <= x"ff740ef1";
		wait for Clk_period;
		Addr <=  "0001110110010";
		Trees_din <= x"09004508";
		wait for Clk_period;
		Addr <=  "0001110110011";
		Trees_din <= x"00fc9804";
		wait for Clk_period;
		Addr <=  "0001110110100";
		Trees_din <= x"002c0ef1";
		wait for Clk_period;
		Addr <=  "0001110110101";
		Trees_din <= x"00980ef1";
		wait for Clk_period;
		Addr <=  "0001110110110";
		Trees_din <= x"0c00c004";
		wait for Clk_period;
		Addr <=  "0001110110111";
		Trees_din <= x"ff7d0ef1";
		wait for Clk_period;
		Addr <=  "0001110111000";
		Trees_din <= x"006f0ef1";
		wait for Clk_period;
		Addr <=  "0001110111001";
		Trees_din <= x"12005904";
		wait for Clk_period;
		Addr <=  "0001110111010";
		Trees_din <= x"00a10ef1";
		wait for Clk_period;
		Addr <=  "0001110111011";
		Trees_din <= x"ffb10ef1";
		wait for Clk_period;
		Addr <=  "0001110111100";
		Trees_din <= x"060c1754";
		wait for Clk_period;
		Addr <=  "0001110111101";
		Trees_din <= x"06013014";
		wait for Clk_period;
		Addr <=  "0001110111110";
		Trees_din <= x"1300ce08";
		wait for Clk_period;
		Addr <=  "0001110111111";
		Trees_din <= x"09004d04";
		wait for Clk_period;
		Addr <=  "0001111000000";
		Trees_din <= x"ff6a101d";
		wait for Clk_period;
		Addr <=  "0001111000001";
		Trees_din <= x"0041101d";
		wait for Clk_period;
		Addr <=  "0001111000010";
		Trees_din <= x"01fddd08";
		wait for Clk_period;
		Addr <=  "0001111000011";
		Trees_din <= x"02fb7804";
		wait for Clk_period;
		Addr <=  "0001111000100";
		Trees_din <= x"000d101d";
		wait for Clk_period;
		Addr <=  "0001111000101";
		Trees_din <= x"00ba101d";
		wait for Clk_period;
		Addr <=  "0001111000110";
		Trees_din <= x"ff8c101d";
		wait for Clk_period;
		Addr <=  "0001111000111";
		Trees_din <= x"1703e520";
		wait for Clk_period;
		Addr <=  "0001111001000";
		Trees_din <= x"1703d010";
		wait for Clk_period;
		Addr <=  "0001111001001";
		Trees_din <= x"15f71808";
		wait for Clk_period;
		Addr <=  "0001111001010";
		Trees_din <= x"07001604";
		wait for Clk_period;
		Addr <=  "0001111001011";
		Trees_din <= x"ff17101d";
		wait for Clk_period;
		Addr <=  "0001111001100";
		Trees_din <= x"0054101d";
		wait for Clk_period;
		Addr <=  "0001111001101";
		Trees_din <= x"11000004";
		wait for Clk_period;
		Addr <=  "0001111001110";
		Trees_din <= x"ffbf101d";
		wait for Clk_period;
		Addr <=  "0001111001111";
		Trees_din <= x"001d101d";
		wait for Clk_period;
		Addr <=  "0001111010000";
		Trees_din <= x"00fd4808";
		wait for Clk_period;
		Addr <=  "0001111010001";
		Trees_din <= x"060af404";
		wait for Clk_period;
		Addr <=  "0001111010010";
		Trees_din <= x"ff3e101d";
		wait for Clk_period;
		Addr <=  "0001111010011";
		Trees_din <= x"0076101d";
		wait for Clk_period;
		Addr <=  "0001111010100";
		Trees_din <= x"05fe4704";
		wait for Clk_period;
		Addr <=  "0001111010101";
		Trees_din <= x"0020101d";
		wait for Clk_period;
		Addr <=  "0001111010110";
		Trees_din <= x"ffa2101d";
		wait for Clk_period;
		Addr <=  "0001111010111";
		Trees_din <= x"1703ec10";
		wait for Clk_period;
		Addr <=  "0001111011000";
		Trees_din <= x"0b00d008";
		wait for Clk_period;
		Addr <=  "0001111011001";
		Trees_din <= x"03fbe904";
		wait for Clk_period;
		Addr <=  "0001111011010";
		Trees_din <= x"ff7f101d";
		wait for Clk_period;
		Addr <=  "0001111011011";
		Trees_din <= x"0057101d";
		wait for Clk_period;
		Addr <=  "0001111011100";
		Trees_din <= x"06060104";
		wait for Clk_period;
		Addr <=  "0001111011101";
		Trees_din <= x"ff9a101d";
		wait for Clk_period;
		Addr <=  "0001111011110";
		Trees_din <= x"00d6101d";
		wait for Clk_period;
		Addr <=  "0001111011111";
		Trees_din <= x"01feff08";
		wait for Clk_period;
		Addr <=  "0001111100000";
		Trees_din <= x"14004a04";
		wait for Clk_period;
		Addr <=  "0001111100001";
		Trees_din <= x"0007101d";
		wait for Clk_period;
		Addr <=  "0001111100010";
		Trees_din <= x"0052101d";
		wait for Clk_period;
		Addr <=  "0001111100011";
		Trees_din <= x"01ff7704";
		wait for Clk_period;
		Addr <=  "0001111100100";
		Trees_din <= x"00c1101d";
		wait for Clk_period;
		Addr <=  "0001111100101";
		Trees_din <= x"0020101d";
		wait for Clk_period;
		Addr <=  "0001111100110";
		Trees_din <= x"10000218";
		wait for Clk_period;
		Addr <=  "0001111100111";
		Trees_din <= x"060d0810";
		wait for Clk_period;
		Addr <=  "0001111101000";
		Trees_din <= x"00fd3404";
		wait for Clk_period;
		Addr <=  "0001111101001";
		Trees_din <= x"fee4101d";
		wait for Clk_period;
		Addr <=  "0001111101010";
		Trees_din <= x"12005508";
		wait for Clk_period;
		Addr <=  "0001111101011";
		Trees_din <= x"03fe1304";
		wait for Clk_period;
		Addr <=  "0001111101100";
		Trees_din <= x"ff7d101d";
		wait for Clk_period;
		Addr <=  "0001111101101";
		Trees_din <= x"fff4101d";
		wait for Clk_period;
		Addr <=  "0001111101110";
		Trees_din <= x"006d101d";
		wait for Clk_period;
		Addr <=  "0001111101111";
		Trees_din <= x"08005004";
		wait for Clk_period;
		Addr <=  "0001111110000";
		Trees_din <= x"0088101d";
		wait for Clk_period;
		Addr <=  "0001111110001";
		Trees_din <= x"ffe5101d";
		wait for Clk_period;
		Addr <=  "0001111110010";
		Trees_din <= x"03028a14";
		wait for Clk_period;
		Addr <=  "0001111110011";
		Trees_din <= x"04066f10";
		wait for Clk_period;
		Addr <=  "0001111110100";
		Trees_din <= x"0b010408";
		wait for Clk_period;
		Addr <=  "0001111110101";
		Trees_din <= x"1e028404";
		wait for Clk_period;
		Addr <=  "0001111110110";
		Trees_din <= x"0096101d";
		wait for Clk_period;
		Addr <=  "0001111110111";
		Trees_din <= x"002d101d";
		wait for Clk_period;
		Addr <=  "0001111111000";
		Trees_din <= x"05fe7804";
		wait for Clk_period;
		Addr <=  "0001111111001";
		Trees_din <= x"ff51101d";
		wait for Clk_period;
		Addr <=  "0001111111010";
		Trees_din <= x"0078101d";
		wait for Clk_period;
		Addr <=  "0001111111011";
		Trees_din <= x"ffb8101d";
		wait for Clk_period;
		Addr <=  "0001111111100";
		Trees_din <= x"1e026108";
		wait for Clk_period;
		Addr <=  "0001111111101";
		Trees_din <= x"00fedc04";
		wait for Clk_period;
		Addr <=  "0001111111110";
		Trees_din <= x"00a1101d";
		wait for Clk_period;
		Addr <=  "0001111111111";
		Trees_din <= x"0024101d";
		wait for Clk_period;
		Addr <=  "0010000000000";
		Trees_din <= x"060e7708";
		wait for Clk_period;
		Addr <=  "0010000000001";
		Trees_din <= x"0f007b04";
		wait for Clk_period;
		Addr <=  "0010000000010";
		Trees_din <= x"002a101d";
		wait for Clk_period;
		Addr <=  "0010000000011";
		Trees_din <= x"ff9b101d";
		wait for Clk_period;
		Addr <=  "0010000000100";
		Trees_din <= x"10001204";
		wait for Clk_period;
		Addr <=  "0010000000101";
		Trees_din <= x"ffc9101d";
		wait for Clk_period;
		Addr <=  "0010000000110";
		Trees_din <= x"007c101d";
		wait for Clk_period;
		Addr <=  "0010000000111";
		Trees_din <= x"060d3258";
		wait for Clk_period;
		Addr <=  "0010000001000";
		Trees_din <= x"06040e28";
		wait for Clk_period;
		Addr <=  "0010000001001";
		Trees_din <= x"0e002f10";
		wait for Clk_period;
		Addr <=  "0010000001010";
		Trees_din <= x"01fd2a08";
		wait for Clk_period;
		Addr <=  "0010000001011";
		Trees_din <= x"0407b704";
		wait for Clk_period;
		Addr <=  "0010000001100";
		Trees_din <= x"ff881129";
		wait for Clk_period;
		Addr <=  "0010000001101";
		Trees_din <= x"00a81129";
		wait for Clk_period;
		Addr <=  "0010000001110";
		Trees_din <= x"0c029604";
		wait for Clk_period;
		Addr <=  "0010000001111";
		Trees_din <= x"ff6c1129";
		wait for Clk_period;
		Addr <=  "0010000010000";
		Trees_din <= x"00021129";
		wait for Clk_period;
		Addr <=  "0010000010001";
		Trees_din <= x"06005808";
		wait for Clk_period;
		Addr <=  "0010000010010";
		Trees_din <= x"1800a704";
		wait for Clk_period;
		Addr <=  "0010000010011";
		Trees_din <= x"ff741129";
		wait for Clk_period;
		Addr <=  "0010000010100";
		Trees_din <= x"00351129";
		wait for Clk_period;
		Addr <=  "0010000010101";
		Trees_din <= x"14004108";
		wait for Clk_period;
		Addr <=  "0010000010110";
		Trees_din <= x"00fe7304";
		wait for Clk_period;
		Addr <=  "0010000010111";
		Trees_din <= x"ff861129";
		wait for Clk_period;
		Addr <=  "0010000011000";
		Trees_din <= x"00a41129";
		wait for Clk_period;
		Addr <=  "0010000011001";
		Trees_din <= x"0d007f04";
		wait for Clk_period;
		Addr <=  "0010000011010";
		Trees_din <= x"ff9b1129";
		wait for Clk_period;
		Addr <=  "0010000011011";
		Trees_din <= x"004d1129";
		wait for Clk_period;
		Addr <=  "0010000011100";
		Trees_din <= x"14005720";
		wait for Clk_period;
		Addr <=  "0010000011101";
		Trees_din <= x"0609e510";
		wait for Clk_period;
		Addr <=  "0010000011110";
		Trees_din <= x"0f007f08";
		wait for Clk_period;
		Addr <=  "0010000011111";
		Trees_din <= x"08004504";
		wait for Clk_period;
		Addr <=  "0010000100000";
		Trees_din <= x"00151129";
		wait for Clk_period;
		Addr <=  "0010000100001";
		Trees_din <= x"ffe41129";
		wait for Clk_period;
		Addr <=  "0010000100010";
		Trees_din <= x"01fc7404";
		wait for Clk_period;
		Addr <=  "0010000100011";
		Trees_din <= x"ffa41129";
		wait for Clk_period;
		Addr <=  "0010000100100";
		Trees_din <= x"00331129";
		wait for Clk_period;
		Addr <=  "0010000100101";
		Trees_din <= x"0f005008";
		wait for Clk_period;
		Addr <=  "0010000100110";
		Trees_din <= x"00fe5a04";
		wait for Clk_period;
		Addr <=  "0010000100111";
		Trees_din <= x"ff2b1129";
		wait for Clk_period;
		Addr <=  "0010000101000";
		Trees_din <= x"00551129";
		wait for Clk_period;
		Addr <=  "0010000101001";
		Trees_din <= x"21000104";
		wait for Clk_period;
		Addr <=  "0010000101010";
		Trees_din <= x"00251129";
		wait for Clk_period;
		Addr <=  "0010000101011";
		Trees_din <= x"00a61129";
		wait for Clk_period;
		Addr <=  "0010000101100";
		Trees_din <= x"0b006f04";
		wait for Clk_period;
		Addr <=  "0010000101101";
		Trees_din <= x"ffe51129";
		wait for Clk_period;
		Addr <=  "0010000101110";
		Trees_din <= x"0c029e08";
		wait for Clk_period;
		Addr <=  "0010000101111";
		Trees_din <= x"0c000004";
		wait for Clk_period;
		Addr <=  "0010000110000";
		Trees_din <= x"003e1129";
		wait for Clk_period;
		Addr <=  "0010000110001";
		Trees_din <= x"00df1129";
		wait for Clk_period;
		Addr <=  "0010000110010";
		Trees_din <= x"fffe1129";
		wait for Clk_period;
		Addr <=  "0010000110011";
		Trees_din <= x"0305bc18";
		wait for Clk_period;
		Addr <=  "0010000110100";
		Trees_din <= x"0f005d08";
		wait for Clk_period;
		Addr <=  "0010000110101";
		Trees_din <= x"09003d04";
		wait for Clk_period;
		Addr <=  "0010000110110";
		Trees_din <= x"00701129";
		wait for Clk_period;
		Addr <=  "0010000110111";
		Trees_din <= x"ff451129";
		wait for Clk_period;
		Addr <=  "0010000111000";
		Trees_din <= x"1ffd1c04";
		wait for Clk_period;
		Addr <=  "0010000111001";
		Trees_din <= x"ffd21129";
		wait for Clk_period;
		Addr <=  "0010000111010";
		Trees_din <= x"0b010a08";
		wait for Clk_period;
		Addr <=  "0010000111011";
		Trees_din <= x"05063404";
		wait for Clk_period;
		Addr <=  "0010000111100";
		Trees_din <= x"00a01129";
		wait for Clk_period;
		Addr <=  "0010000111101";
		Trees_din <= x"00331129";
		wait for Clk_period;
		Addr <=  "0010000111110";
		Trees_din <= x"00011129";
		wait for Clk_period;
		Addr <=  "0010000111111";
		Trees_din <= x"01fc3108";
		wait for Clk_period;
		Addr <=  "0010001000000";
		Trees_din <= x"0e002504";
		wait for Clk_period;
		Addr <=  "0010001000001";
		Trees_din <= x"ff511129";
		wait for Clk_period;
		Addr <=  "0010001000010";
		Trees_din <= x"003f1129";
		wait for Clk_period;
		Addr <=  "0010001000011";
		Trees_din <= x"0309a404";
		wait for Clk_period;
		Addr <=  "0010001000100";
		Trees_din <= x"00931129";
		wait for Clk_period;
		Addr <=  "0010001000101";
		Trees_din <= x"0d006a04";
		wait for Clk_period;
		Addr <=  "0010001000110";
		Trees_din <= x"00551129";
		wait for Clk_period;
		Addr <=  "0010001000111";
		Trees_din <= x"1afbf104";
		wait for Clk_period;
		Addr <=  "0010001001000";
		Trees_din <= x"ff761129";
		wait for Clk_period;
		Addr <=  "0010001001001";
		Trees_din <= x"002d1129";
		wait for Clk_period;
		Addr <=  "0010001001010";
		Trees_din <= x"060d6854";
		wait for Clk_period;
		Addr <=  "0010001001011";
		Trees_din <= x"06013014";
		wait for Clk_period;
		Addr <=  "0010001001100";
		Trees_din <= x"1300ce08";
		wait for Clk_period;
		Addr <=  "0010001001101";
		Trees_din <= x"09004d04";
		wait for Clk_period;
		Addr <=  "0010001001110";
		Trees_din <= x"ff6d121d";
		wait for Clk_period;
		Addr <=  "0010001001111";
		Trees_din <= x"003e121d";
		wait for Clk_period;
		Addr <=  "0010001010000";
		Trees_din <= x"0f008508";
		wait for Clk_period;
		Addr <=  "0010001010001";
		Trees_din <= x"1703b004";
		wait for Clk_period;
		Addr <=  "0010001010010";
		Trees_din <= x"00b0121d";
		wait for Clk_period;
		Addr <=  "0010001010011";
		Trees_din <= x"000f121d";
		wait for Clk_period;
		Addr <=  "0010001010100";
		Trees_din <= x"ff95121d";
		wait for Clk_period;
		Addr <=  "0010001010101";
		Trees_din <= x"1f028420";
		wait for Clk_period;
		Addr <=  "0010001010110";
		Trees_din <= x"1b028310";
		wait for Clk_period;
		Addr <=  "0010001010111";
		Trees_din <= x"14004708";
		wait for Clk_period;
		Addr <=  "0010001011000";
		Trees_din <= x"09004d04";
		wait for Clk_period;
		Addr <=  "0010001011001";
		Trees_din <= x"000d121d";
		wait for Clk_period;
		Addr <=  "0010001011010";
		Trees_din <= x"ff7b121d";
		wait for Clk_period;
		Addr <=  "0010001011011";
		Trees_din <= x"1c025404";
		wait for Clk_period;
		Addr <=  "0010001011100";
		Trees_din <= x"ffff121d";
		wait for Clk_period;
		Addr <=  "0010001011101";
		Trees_din <= x"0049121d";
		wait for Clk_period;
		Addr <=  "0010001011110";
		Trees_din <= x"0406d408";
		wait for Clk_period;
		Addr <=  "0010001011111";
		Trees_din <= x"08005b04";
		wait for Clk_period;
		Addr <=  "0010001100000";
		Trees_din <= x"008e121d";
		wait for Clk_period;
		Addr <=  "0010001100001";
		Trees_din <= x"ff99121d";
		wait for Clk_period;
		Addr <=  "0010001100010";
		Trees_din <= x"05fc5204";
		wait for Clk_period;
		Addr <=  "0010001100011";
		Trees_din <= x"0063121d";
		wait for Clk_period;
		Addr <=  "0010001100100";
		Trees_din <= x"ff76121d";
		wait for Clk_period;
		Addr <=  "0010001100101";
		Trees_din <= x"12003c10";
		wait for Clk_period;
		Addr <=  "0010001100110";
		Trees_din <= x"1001ca08";
		wait for Clk_period;
		Addr <=  "0010001100111";
		Trees_din <= x"01fd8704";
		wait for Clk_period;
		Addr <=  "0010001101000";
		Trees_din <= x"ff6e121d";
		wait for Clk_period;
		Addr <=  "0010001101001";
		Trees_din <= x"003d121d";
		wait for Clk_period;
		Addr <=  "0010001101010";
		Trees_din <= x"1300ba04";
		wait for Clk_period;
		Addr <=  "0010001101011";
		Trees_din <= x"0062121d";
		wait for Clk_period;
		Addr <=  "0010001101100";
		Trees_din <= x"ff0c121d";
		wait for Clk_period;
		Addr <=  "0010001101101";
		Trees_din <= x"0c030108";
		wait for Clk_period;
		Addr <=  "0010001101110";
		Trees_din <= x"12004a04";
		wait for Clk_period;
		Addr <=  "0010001101111";
		Trees_din <= x"0045121d";
		wait for Clk_period;
		Addr <=  "0010001110000";
		Trees_din <= x"ffd4121d";
		wait for Clk_period;
		Addr <=  "0010001110001";
		Trees_din <= x"13009904";
		wait for Clk_period;
		Addr <=  "0010001110010";
		Trees_din <= x"00aa121d";
		wait for Clk_period;
		Addr <=  "0010001110011";
		Trees_din <= x"ff74121d";
		wait for Clk_period;
		Addr <=  "0010001110100";
		Trees_din <= x"03036808";
		wait for Clk_period;
		Addr <=  "0010001110101";
		Trees_din <= x"1102ac04";
		wait for Clk_period;
		Addr <=  "0010001110110";
		Trees_din <= x"009b121d";
		wait for Clk_period;
		Addr <=  "0010001110111";
		Trees_din <= x"fffe121d";
		wait for Clk_period;
		Addr <=  "0010001111000";
		Trees_din <= x"2004000c";
		wait for Clk_period;
		Addr <=  "0010001111001";
		Trees_din <= x"0d009808";
		wait for Clk_period;
		Addr <=  "0010001111010";
		Trees_din <= x"0a004604";
		wait for Clk_period;
		Addr <=  "0010001111011";
		Trees_din <= x"ff5a121d";
		wait for Clk_period;
		Addr <=  "0010001111100";
		Trees_din <= x"0029121d";
		wait for Clk_period;
		Addr <=  "0010001111101";
		Trees_din <= x"005c121d";
		wait for Clk_period;
		Addr <=  "0010001111110";
		Trees_din <= x"04f9fd10";
		wait for Clk_period;
		Addr <=  "0010001111111";
		Trees_din <= x"08004208";
		wait for Clk_period;
		Addr <=  "0010010000000";
		Trees_din <= x"07faca04";
		wait for Clk_period;
		Addr <=  "0010010000001";
		Trees_din <= x"ff74121d";
		wait for Clk_period;
		Addr <=  "0010010000010";
		Trees_din <= x"005d121d";
		wait for Clk_period;
		Addr <=  "0010010000011";
		Trees_din <= x"0501c304";
		wait for Clk_period;
		Addr <=  "0010010000100";
		Trees_din <= x"001e121d";
		wait for Clk_period;
		Addr <=  "0010010000101";
		Trees_din <= x"007a121d";
		wait for Clk_period;
		Addr <=  "0010010000110";
		Trees_din <= x"0097121d";
		wait for Clk_period;
		Addr <=  "0010010000111";
		Trees_din <= x"060d6830";
		wait for Clk_period;
		Addr <=  "0010010001000";
		Trees_din <= x"0002622c";
		wait for Clk_period;
		Addr <=  "0010010001001";
		Trees_din <= x"14005718";
		wait for Clk_period;
		Addr <=  "0010010001010";
		Trees_din <= x"06ffb808";
		wait for Clk_period;
		Addr <=  "0010010001011";
		Trees_din <= x"0c029604";
		wait for Clk_period;
		Addr <=  "0010010001100";
		Trees_din <= x"ff7812c9";
		wait for Clk_period;
		Addr <=  "0010010001101";
		Trees_din <= x"002012c9";
		wait for Clk_period;
		Addr <=  "0010010001110";
		Trees_din <= x"03fa3e08";
		wait for Clk_period;
		Addr <=  "0010010001111";
		Trees_din <= x"1300dc04";
		wait for Clk_period;
		Addr <=  "0010010010000";
		Trees_din <= x"006c12c9";
		wait for Clk_period;
		Addr <=  "0010010010001";
		Trees_din <= x"ff5912c9";
		wait for Clk_period;
		Addr <=  "0010010010010";
		Trees_din <= x"03fabd04";
		wait for Clk_period;
		Addr <=  "0010010010011";
		Trees_din <= x"ffcc12c9";
		wait for Clk_period;
		Addr <=  "0010010010100";
		Trees_din <= x"000f12c9";
		wait for Clk_period;
		Addr <=  "0010010010101";
		Trees_din <= x"12005c04";
		wait for Clk_period;
		Addr <=  "0010010010110";
		Trees_din <= x"ffbe12c9";
		wait for Clk_period;
		Addr <=  "0010010010111";
		Trees_din <= x"02fa4d08";
		wait for Clk_period;
		Addr <=  "0010010011000";
		Trees_din <= x"08004e04";
		wait for Clk_period;
		Addr <=  "0010010011001";
		Trees_din <= x"ff8612c9";
		wait for Clk_period;
		Addr <=  "0010010011010";
		Trees_din <= x"007812c9";
		wait for Clk_period;
		Addr <=  "0010010011011";
		Trees_din <= x"12006104";
		wait for Clk_period;
		Addr <=  "0010010011100";
		Trees_din <= x"00d312c9";
		wait for Clk_period;
		Addr <=  "0010010011101";
		Trees_din <= x"004612c9";
		wait for Clk_period;
		Addr <=  "0010010011110";
		Trees_din <= x"ff7512c9";
		wait for Clk_period;
		Addr <=  "0010010011111";
		Trees_din <= x"03028a04";
		wait for Clk_period;
		Addr <=  "0010010100000";
		Trees_din <= x"009712c9";
		wait for Clk_period;
		Addr <=  "0010010100001";
		Trees_din <= x"20040010";
		wait for Clk_period;
		Addr <=  "0010010100010";
		Trees_din <= x"060f690c";
		wait for Clk_period;
		Addr <=  "0010010100011";
		Trees_din <= x"14003a04";
		wait for Clk_period;
		Addr <=  "0010010100100";
		Trees_din <= x"002712c9";
		wait for Clk_period;
		Addr <=  "0010010100101";
		Trees_din <= x"0a000b04";
		wait for Clk_period;
		Addr <=  "0010010100110";
		Trees_din <= x"ff5c12c9";
		wait for Clk_period;
		Addr <=  "0010010100111";
		Trees_din <= x"ffdc12c9";
		wait for Clk_period;
		Addr <=  "0010010101000";
		Trees_din <= x"005b12c9";
		wait for Clk_period;
		Addr <=  "0010010101001";
		Trees_din <= x"0a01760c";
		wait for Clk_period;
		Addr <=  "0010010101010";
		Trees_din <= x"0b00ea04";
		wait for Clk_period;
		Addr <=  "0010010101011";
		Trees_din <= x"009012c9";
		wait for Clk_period;
		Addr <=  "0010010101100";
		Trees_din <= x"02fe3f04";
		wait for Clk_period;
		Addr <=  "0010010101101";
		Trees_din <= x"005b12c9";
		wait for Clk_period;
		Addr <=  "0010010101110";
		Trees_din <= x"ffbc12c9";
		wait for Clk_period;
		Addr <=  "0010010101111";
		Trees_din <= x"1b027004";
		wait for Clk_period;
		Addr <=  "0010010110000";
		Trees_din <= x"ffa612c9";
		wait for Clk_period;
		Addr <=  "0010010110001";
		Trees_din <= x"005a12c9";
		wait for Clk_period;
		Addr <=  "0010010110010";
		Trees_din <= x"060d6838";
		wait for Clk_period;
		Addr <=  "0010010110011";
		Trees_din <= x"00026234";
		wait for Clk_period;
		Addr <=  "0010010110100";
		Trees_din <= x"14005720";
		wait for Clk_period;
		Addr <=  "0010010110101";
		Trees_din <= x"06013010";
		wait for Clk_period;
		Addr <=  "0010010110110";
		Trees_din <= x"1300ce08";
		wait for Clk_period;
		Addr <=  "0010010110111";
		Trees_din <= x"0a000004";
		wait for Clk_period;
		Addr <=  "0010010111000";
		Trees_din <= x"fff1138d";
		wait for Clk_period;
		Addr <=  "0010010111001";
		Trees_din <= x"ff75138d";
		wait for Clk_period;
		Addr <=  "0010010111010";
		Trees_din <= x"01fddd04";
		wait for Clk_period;
		Addr <=  "0010010111011";
		Trees_din <= x"0084138d";
		wait for Clk_period;
		Addr <=  "0010010111100";
		Trees_din <= x"ffad138d";
		wait for Clk_period;
		Addr <=  "0010010111101";
		Trees_din <= x"1f028408";
		wait for Clk_period;
		Addr <=  "0010010111110";
		Trees_din <= x"1b028304";
		wait for Clk_period;
		Addr <=  "0010010111111";
		Trees_din <= x"000c138d";
		wait for Clk_period;
		Addr <=  "0010011000000";
		Trees_din <= x"0059138d";
		wait for Clk_period;
		Addr <=  "0010011000001";
		Trees_din <= x"03fcaa04";
		wait for Clk_period;
		Addr <=  "0010011000010";
		Trees_din <= x"ffbc138d";
		wait for Clk_period;
		Addr <=  "0010011000011";
		Trees_din <= x"0014138d";
		wait for Clk_period;
		Addr <=  "0010011000100";
		Trees_din <= x"0405c504";
		wait for Clk_period;
		Addr <=  "0010011000101";
		Trees_din <= x"00a5138d";
		wait for Clk_period;
		Addr <=  "0010011000110";
		Trees_din <= x"05fd7208";
		wait for Clk_period;
		Addr <=  "0010011000111";
		Trees_din <= x"0a000004";
		wait for Clk_period;
		Addr <=  "0010011001000";
		Trees_din <= x"ffdd138d";
		wait for Clk_period;
		Addr <=  "0010011001001";
		Trees_din <= x"ff83138d";
		wait for Clk_period;
		Addr <=  "0010011001010";
		Trees_din <= x"0b008f04";
		wait for Clk_period;
		Addr <=  "0010011001011";
		Trees_din <= x"00bc138d";
		wait for Clk_period;
		Addr <=  "0010011001100";
		Trees_din <= x"ffe7138d";
		wait for Clk_period;
		Addr <=  "0010011001101";
		Trees_din <= x"ff7a138d";
		wait for Clk_period;
		Addr <=  "0010011001110";
		Trees_din <= x"03028a04";
		wait for Clk_period;
		Addr <=  "0010011001111";
		Trees_din <= x"0094138d";
		wait for Clk_period;
		Addr <=  "0010011010000";
		Trees_din <= x"20040010";
		wait for Clk_period;
		Addr <=  "0010011010001";
		Trees_din <= x"060f690c";
		wait for Clk_period;
		Addr <=  "0010011010010";
		Trees_din <= x"08004404";
		wait for Clk_period;
		Addr <=  "0010011010011";
		Trees_din <= x"0024138d";
		wait for Clk_period;
		Addr <=  "0010011010100";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "0010011010101";
		Trees_din <= x"ffd4138d";
		wait for Clk_period;
		Addr <=  "0010011010110";
		Trees_din <= x"ff6d138d";
		wait for Clk_period;
		Addr <=  "0010011010111";
		Trees_din <= x"0056138d";
		wait for Clk_period;
		Addr <=  "0010011011000";
		Trees_din <= x"0f008710";
		wait for Clk_period;
		Addr <=  "0010011011001";
		Trees_din <= x"0b00ea08";
		wait for Clk_period;
		Addr <=  "0010011011010";
		Trees_din <= x"17023104";
		wait for Clk_period;
		Addr <=  "0010011011011";
		Trees_din <= x"0014138d";
		wait for Clk_period;
		Addr <=  "0010011011100";
		Trees_din <= x"008c138d";
		wait for Clk_period;
		Addr <=  "0010011011101";
		Trees_din <= x"02fe3f04";
		wait for Clk_period;
		Addr <=  "0010011011110";
		Trees_din <= x"0054138d";
		wait for Clk_period;
		Addr <=  "0010011011111";
		Trees_din <= x"ffc1138d";
		wait for Clk_period;
		Addr <=  "0010011100000";
		Trees_din <= x"05025504";
		wait for Clk_period;
		Addr <=  "0010011100001";
		Trees_din <= x"003b138d";
		wait for Clk_period;
		Addr <=  "0010011100010";
		Trees_din <= x"ffab138d";
		wait for Clk_period;
		Addr <=  "0010011100011";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0010011100100";
		Trees_din <= x"060d6844";
		wait for Clk_period;
		Addr <=  "0010011100101";
		Trees_din <= x"00026240";
		wait for Clk_period;
		Addr <=  "0010011100110";
		Trees_din <= x"00fd9420";
		wait for Clk_period;
		Addr <=  "0010011100111";
		Trees_din <= x"15f99810";
		wait for Clk_period;
		Addr <=  "0010011101000";
		Trees_din <= x"1afa5308";
		wait for Clk_period;
		Addr <=  "0010011101001";
		Trees_din <= x"07fe0a04";
		wait for Clk_period;
		Addr <=  "0010011101010";
		Trees_din <= x"007c1455";
		wait for Clk_period;
		Addr <=  "0010011101011";
		Trees_din <= x"fec11455";
		wait for Clk_period;
		Addr <=  "0010011101100";
		Trees_din <= x"0c031404";
		wait for Clk_period;
		Addr <=  "0010011101101";
		Trees_din <= x"ffed1455";
		wait for Clk_period;
		Addr <=  "0010011101110";
		Trees_din <= x"007f1455";
		wait for Clk_period;
		Addr <=  "0010011101111";
		Trees_din <= x"05fec608";
		wait for Clk_period;
		Addr <=  "0010011110000";
		Trees_din <= x"08004f04";
		wait for Clk_period;
		Addr <=  "0010011110001";
		Trees_din <= x"00881455";
		wait for Clk_period;
		Addr <=  "0010011110010";
		Trees_din <= x"ffe61455";
		wait for Clk_period;
		Addr <=  "0010011110011";
		Trees_din <= x"0e002c04";
		wait for Clk_period;
		Addr <=  "0010011110100";
		Trees_din <= x"ff451455";
		wait for Clk_period;
		Addr <=  "0010011110101";
		Trees_din <= x"005b1455";
		wait for Clk_period;
		Addr <=  "0010011110110";
		Trees_din <= x"0c02b610";
		wait for Clk_period;
		Addr <=  "0010011110111";
		Trees_din <= x"1002d508";
		wait for Clk_period;
		Addr <=  "0010011111000";
		Trees_din <= x"17029704";
		wait for Clk_period;
		Addr <=  "0010011111001";
		Trees_din <= x"005a1455";
		wait for Clk_period;
		Addr <=  "0010011111010";
		Trees_din <= x"00121455";
		wait for Clk_period;
		Addr <=  "0010011111011";
		Trees_din <= x"0e003d04";
		wait for Clk_period;
		Addr <=  "0010011111100";
		Trees_din <= x"ffa01455";
		wait for Clk_period;
		Addr <=  "0010011111101";
		Trees_din <= x"00391455";
		wait for Clk_period;
		Addr <=  "0010011111110";
		Trees_din <= x"0f007108";
		wait for Clk_period;
		Addr <=  "0010011111111";
		Trees_din <= x"03fbd904";
		wait for Clk_period;
		Addr <=  "0010100000000";
		Trees_din <= x"00f01455";
		wait for Clk_period;
		Addr <=  "0010100000001";
		Trees_din <= x"00061455";
		wait for Clk_period;
		Addr <=  "0010100000010";
		Trees_din <= x"0f008c04";
		wait for Clk_period;
		Addr <=  "0010100000011";
		Trees_din <= x"ffa41455";
		wait for Clk_period;
		Addr <=  "0010100000100";
		Trees_din <= x"006d1455";
		wait for Clk_period;
		Addr <=  "0010100000101";
		Trees_din <= x"ff811455";
		wait for Clk_period;
		Addr <=  "0010100000110";
		Trees_din <= x"03028a04";
		wait for Clk_period;
		Addr <=  "0010100000111";
		Trees_din <= x"00911455";
		wait for Clk_period;
		Addr <=  "0010100001000";
		Trees_din <= x"2004000c";
		wait for Clk_period;
		Addr <=  "0010100001001";
		Trees_din <= x"00fdd608";
		wait for Clk_period;
		Addr <=  "0010100001010";
		Trees_din <= x"09003f04";
		wait for Clk_period;
		Addr <=  "0010100001011";
		Trees_din <= x"001c1455";
		wait for Clk_period;
		Addr <=  "0010100001100";
		Trees_din <= x"ff7b1455";
		wait for Clk_period;
		Addr <=  "0010100001101";
		Trees_din <= x"00311455";
		wait for Clk_period;
		Addr <=  "0010100001110";
		Trees_din <= x"0a017608";
		wait for Clk_period;
		Addr <=  "0010100001111";
		Trees_din <= x"0b00ea04";
		wait for Clk_period;
		Addr <=  "0010100010000";
		Trees_din <= x"00851455";
		wait for Clk_period;
		Addr <=  "0010100010001";
		Trees_din <= x"000f1455";
		wait for Clk_period;
		Addr <=  "0010100010010";
		Trees_din <= x"0a01a504";
		wait for Clk_period;
		Addr <=  "0010100010011";
		Trees_din <= x"ff9d1455";
		wait for Clk_period;
		Addr <=  "0010100010100";
		Trees_din <= x"00431455";
		wait for Clk_period;
		Addr <=  "0010100010101";
		Trees_din <= x"060d6860";
		wait for Clk_period;
		Addr <=  "0010100010110";
		Trees_din <= x"06040e24";
		wait for Clk_period;
		Addr <=  "0010100010111";
		Trees_din <= x"00fdd608";
		wait for Clk_period;
		Addr <=  "0010100011000";
		Trees_din <= x"22000204";
		wait for Clk_period;
		Addr <=  "0010100011001";
		Trees_din <= x"ff751551";
		wait for Clk_period;
		Addr <=  "0010100011010";
		Trees_din <= x"fff11551";
		wait for Clk_period;
		Addr <=  "0010100011011";
		Trees_din <= x"0e002f10";
		wait for Clk_period;
		Addr <=  "0010100011100";
		Trees_din <= x"00fea808";
		wait for Clk_period;
		Addr <=  "0010100011101";
		Trees_din <= x"01fd2a04";
		wait for Clk_period;
		Addr <=  "0010100011110";
		Trees_din <= x"00c41551";
		wait for Clk_period;
		Addr <=  "0010100011111";
		Trees_din <= x"ff9f1551";
		wait for Clk_period;
		Addr <=  "0010100100000";
		Trees_din <= x"0c028804";
		wait for Clk_period;
		Addr <=  "0010100100001";
		Trees_din <= x"ff741551";
		wait for Clk_period;
		Addr <=  "0010100100010";
		Trees_din <= x"00161551";
		wait for Clk_period;
		Addr <=  "0010100100011";
		Trees_din <= x"05fc0504";
		wait for Clk_period;
		Addr <=  "0010100100100";
		Trees_din <= x"ff821551";
		wait for Clk_period;
		Addr <=  "0010100100101";
		Trees_din <= x"05fc3104";
		wait for Clk_period;
		Addr <=  "0010100100110";
		Trees_din <= x"00c11551";
		wait for Clk_period;
		Addr <=  "0010100100111";
		Trees_din <= x"00091551";
		wait for Clk_period;
		Addr <=  "0010100101000";
		Trees_din <= x"01fd9920";
		wait for Clk_period;
		Addr <=  "0010100101001";
		Trees_din <= x"1300aa10";
		wait for Clk_period;
		Addr <=  "0010100101010";
		Trees_din <= x"03fbdf08";
		wait for Clk_period;
		Addr <=  "0010100101011";
		Trees_din <= x"0607cf04";
		wait for Clk_period;
		Addr <=  "0010100101100";
		Trees_din <= x"00011551";
		wait for Clk_period;
		Addr <=  "0010100101101";
		Trees_din <= x"ff681551";
		wait for Clk_period;
		Addr <=  "0010100101110";
		Trees_din <= x"09004704";
		wait for Clk_period;
		Addr <=  "0010100101111";
		Trees_din <= x"ffea1551";
		wait for Clk_period;
		Addr <=  "0010100110000";
		Trees_din <= x"004d1551";
		wait for Clk_period;
		Addr <=  "0010100110001";
		Trees_din <= x"0d006d08";
		wait for Clk_period;
		Addr <=  "0010100110010";
		Trees_din <= x"1000bf04";
		wait for Clk_period;
		Addr <=  "0010100110011";
		Trees_din <= x"000c1551";
		wait for Clk_period;
		Addr <=  "0010100110100";
		Trees_din <= x"00ad1551";
		wait for Clk_period;
		Addr <=  "0010100110101";
		Trees_din <= x"10033e04";
		wait for Clk_period;
		Addr <=  "0010100110110";
		Trees_din <= x"000b1551";
		wait for Clk_period;
		Addr <=  "0010100110111";
		Trees_din <= x"ff651551";
		wait for Clk_period;
		Addr <=  "0010100111000";
		Trees_din <= x"01fda70c";
		wait for Clk_period;
		Addr <=  "0010100111001";
		Trees_din <= x"1b024704";
		wait for Clk_period;
		Addr <=  "0010100111010";
		Trees_din <= x"ff491551";
		wait for Clk_period;
		Addr <=  "0010100111011";
		Trees_din <= x"18007004";
		wait for Clk_period;
		Addr <=  "0010100111100";
		Trees_din <= x"00de1551";
		wait for Clk_period;
		Addr <=  "0010100111101";
		Trees_din <= x"00291551";
		wait for Clk_period;
		Addr <=  "0010100111110";
		Trees_din <= x"02faf208";
		wait for Clk_period;
		Addr <=  "0010100111111";
		Trees_din <= x"02fa4504";
		wait for Clk_period;
		Addr <=  "0010101000000";
		Trees_din <= x"fffa1551";
		wait for Clk_period;
		Addr <=  "0010101000001";
		Trees_din <= x"00491551";
		wait for Clk_period;
		Addr <=  "0010101000010";
		Trees_din <= x"02faf804";
		wait for Clk_period;
		Addr <=  "0010101000011";
		Trees_din <= x"ff621551";
		wait for Clk_period;
		Addr <=  "0010101000100";
		Trees_din <= x"00041551";
		wait for Clk_period;
		Addr <=  "0010101000101";
		Trees_din <= x"03028a04";
		wait for Clk_period;
		Addr <=  "0010101000110";
		Trees_din <= x"008f1551";
		wait for Clk_period;
		Addr <=  "0010101000111";
		Trees_din <= x"060e9010";
		wait for Clk_period;
		Addr <=  "0010101001000";
		Trees_din <= x"19000c0c";
		wait for Clk_period;
		Addr <=  "0010101001001";
		Trees_din <= x"09004308";
		wait for Clk_period;
		Addr <=  "0010101001010";
		Trees_din <= x"10005a04";
		wait for Clk_period;
		Addr <=  "0010101001011";
		Trees_din <= x"00071551";
		wait for Clk_period;
		Addr <=  "0010101001100";
		Trees_din <= x"ff891551";
		wait for Clk_period;
		Addr <=  "0010101001101";
		Trees_din <= x"00421551";
		wait for Clk_period;
		Addr <=  "0010101001110";
		Trees_din <= x"00581551";
		wait for Clk_period;
		Addr <=  "0010101001111";
		Trees_din <= x"030aad08";
		wait for Clk_period;
		Addr <=  "0010101010000";
		Trees_din <= x"09004504";
		wait for Clk_period;
		Addr <=  "0010101010001";
		Trees_din <= x"00861551";
		wait for Clk_period;
		Addr <=  "0010101010010";
		Trees_din <= x"00131551";
		wait for Clk_period;
		Addr <=  "0010101010011";
		Trees_din <= x"fff21551";
		wait for Clk_period;
		Addr <=  "0010101010100";
		Trees_din <= x"060d687c";
		wait for Clk_period;
		Addr <=  "0010101010101";
		Trees_din <= x"10008a3c";
		wait for Clk_period;
		Addr <=  "0010101010110";
		Trees_din <= x"01fefb20";
		wait for Clk_period;
		Addr <=  "0010101010111";
		Trees_din <= x"11000810";
		wait for Clk_period;
		Addr <=  "0010101011000";
		Trees_din <= x"03fbe408";
		wait for Clk_period;
		Addr <=  "0010101011001";
		Trees_din <= x"02faa604";
		wait for Clk_period;
		Addr <=  "0010101011010";
		Trees_din <= x"0016168d";
		wait for Clk_period;
		Addr <=  "0010101011011";
		Trees_din <= x"ff73168d";
		wait for Clk_period;
		Addr <=  "0010101011100";
		Trees_din <= x"06070104";
		wait for Clk_period;
		Addr <=  "0010101011101";
		Trees_din <= x"ffd2168d";
		wait for Clk_period;
		Addr <=  "0010101011110";
		Trees_din <= x"0019168d";
		wait for Clk_period;
		Addr <=  "0010101011111";
		Trees_din <= x"0c013108";
		wait for Clk_period;
		Addr <=  "0010101100000";
		Trees_din <= x"0c00fe04";
		wait for Clk_period;
		Addr <=  "0010101100001";
		Trees_din <= x"001e168d";
		wait for Clk_period;
		Addr <=  "0010101100010";
		Trees_din <= x"ffa3168d";
		wait for Clk_period;
		Addr <=  "0010101100011";
		Trees_din <= x"0a004504";
		wait for Clk_period;
		Addr <=  "0010101100100";
		Trees_din <= x"0001168d";
		wait for Clk_period;
		Addr <=  "0010101100101";
		Trees_din <= x"0082168d";
		wait for Clk_period;
		Addr <=  "0010101100110";
		Trees_din <= x"01ff7710";
		wait for Clk_period;
		Addr <=  "0010101100111";
		Trees_din <= x"03fe9b08";
		wait for Clk_period;
		Addr <=  "0010101101000";
		Trees_din <= x"02fd1804";
		wait for Clk_period;
		Addr <=  "0010101101001";
		Trees_din <= x"00b6168d";
		wait for Clk_period;
		Addr <=  "0010101101010";
		Trees_din <= x"ffe3168d";
		wait for Clk_period;
		Addr <=  "0010101101011";
		Trees_din <= x"09004304";
		wait for Clk_period;
		Addr <=  "0010101101100";
		Trees_din <= x"0073168d";
		wait for Clk_period;
		Addr <=  "0010101101101";
		Trees_din <= x"ff65168d";
		wait for Clk_period;
		Addr <=  "0010101101110";
		Trees_din <= x"0b00f208";
		wait for Clk_period;
		Addr <=  "0010101101111";
		Trees_din <= x"09003e04";
		wait for Clk_period;
		Addr <=  "0010101110000";
		Trees_din <= x"ff87168d";
		wait for Clk_period;
		Addr <=  "0010101110001";
		Trees_din <= x"003b168d";
		wait for Clk_period;
		Addr <=  "0010101110010";
		Trees_din <= x"0091168d";
		wait for Clk_period;
		Addr <=  "0010101110011";
		Trees_din <= x"1000cd20";
		wait for Clk_period;
		Addr <=  "0010101110100";
		Trees_din <= x"02faea10";
		wait for Clk_period;
		Addr <=  "0010101110101";
		Trees_din <= x"19000208";
		wait for Clk_period;
		Addr <=  "0010101110110";
		Trees_din <= x"00fed804";
		wait for Clk_period;
		Addr <=  "0010101110111";
		Trees_din <= x"ff8b168d";
		wait for Clk_period;
		Addr <=  "0010101111000";
		Trees_din <= x"005c168d";
		wait for Clk_period;
		Addr <=  "0010101111001";
		Trees_din <= x"07003104";
		wait for Clk_period;
		Addr <=  "0010101111010";
		Trees_din <= x"00e6168d";
		wait for Clk_period;
		Addr <=  "0010101111011";
		Trees_din <= x"ff9d168d";
		wait for Clk_period;
		Addr <=  "0010101111100";
		Trees_din <= x"02fb7808";
		wait for Clk_period;
		Addr <=  "0010101111101";
		Trees_din <= x"00feb204";
		wait for Clk_period;
		Addr <=  "0010101111110";
		Trees_din <= x"fee9168d";
		wait for Clk_period;
		Addr <=  "0010101111111";
		Trees_din <= x"fff7168d";
		wait for Clk_period;
		Addr <=  "0010110000000";
		Trees_din <= x"1000c604";
		wait for Clk_period;
		Addr <=  "0010110000001";
		Trees_din <= x"ffda168d";
		wait for Clk_period;
		Addr <=  "0010110000010";
		Trees_din <= x"ff1a168d";
		wait for Clk_period;
		Addr <=  "0010110000011";
		Trees_din <= x"11001410";
		wait for Clk_period;
		Addr <=  "0010110000100";
		Trees_din <= x"1afbdd08";
		wait for Clk_period;
		Addr <=  "0010110000101";
		Trees_din <= x"13009904";
		wait for Clk_period;
		Addr <=  "0010110000110";
		Trees_din <= x"005f168d";
		wait for Clk_period;
		Addr <=  "0010110000111";
		Trees_din <= x"ffbc168d";
		wait for Clk_period;
		Addr <=  "0010110001000";
		Trees_din <= x"07fed204";
		wait for Clk_period;
		Addr <=  "0010110001001";
		Trees_din <= x"0004168d";
		wait for Clk_period;
		Addr <=  "0010110001010";
		Trees_din <= x"00a1168d";
		wait for Clk_period;
		Addr <=  "0010110001011";
		Trees_din <= x"1c027208";
		wait for Clk_period;
		Addr <=  "0010110001100";
		Trees_din <= x"0c010a04";
		wait for Clk_period;
		Addr <=  "0010110001101";
		Trees_din <= x"001d168d";
		wait for Clk_period;
		Addr <=  "0010110001110";
		Trees_din <= x"ffa3168d";
		wait for Clk_period;
		Addr <=  "0010110001111";
		Trees_din <= x"10010104";
		wait for Clk_period;
		Addr <=  "0010110010000";
		Trees_din <= x"005a168d";
		wait for Clk_period;
		Addr <=  "0010110010001";
		Trees_din <= x"fffe168d";
		wait for Clk_period;
		Addr <=  "0010110010010";
		Trees_din <= x"03028a04";
		wait for Clk_period;
		Addr <=  "0010110010011";
		Trees_din <= x"008c168d";
		wait for Clk_period;
		Addr <=  "0010110010100";
		Trees_din <= x"2004000c";
		wait for Clk_period;
		Addr <=  "0010110010101";
		Trees_din <= x"00fdd608";
		wait for Clk_period;
		Addr <=  "0010110010110";
		Trees_din <= x"10005a04";
		wait for Clk_period;
		Addr <=  "0010110010111";
		Trees_din <= x"0000168d";
		wait for Clk_period;
		Addr <=  "0010110011000";
		Trees_din <= x"ff88168d";
		wait for Clk_period;
		Addr <=  "0010110011001";
		Trees_din <= x"0029168d";
		wait for Clk_period;
		Addr <=  "0010110011010";
		Trees_din <= x"04f9fd0c";
		wait for Clk_period;
		Addr <=  "0010110011011";
		Trees_din <= x"08004208";
		wait for Clk_period;
		Addr <=  "0010110011100";
		Trees_din <= x"0c00f704";
		wait for Clk_period;
		Addr <=  "0010110011101";
		Trees_din <= x"ffa3168d";
		wait for Clk_period;
		Addr <=  "0010110011110";
		Trees_din <= x"0001168d";
		wait for Clk_period;
		Addr <=  "0010110011111";
		Trees_din <= x"004c168d";
		wait for Clk_period;
		Addr <=  "0010110100000";
		Trees_din <= x"12004b04";
		wait for Clk_period;
		Addr <=  "0010110100001";
		Trees_din <= x"0084168d";
		wait for Clk_period;
		Addr <=  "0010110100010";
		Trees_din <= x"000b168d";
		wait for Clk_period;
		Addr <=  "0010110100011";
		Trees_din <= x"060d6874";
		wait for Clk_period;
		Addr <=  "0010110100100";
		Trees_din <= x"05fe3938";
		wait for Clk_period;
		Addr <=  "0010110100101";
		Trees_din <= x"03fcf218";
		wait for Clk_period;
		Addr <=  "0010110100110";
		Trees_din <= x"01fc2708";
		wait for Clk_period;
		Addr <=  "0010110100111";
		Trees_din <= x"04041504";
		wait for Clk_period;
		Addr <=  "0010110101000";
		Trees_din <= x"000417b9";
		wait for Clk_period;
		Addr <=  "0010110101001";
		Trees_din <= x"ff3b17b9";
		wait for Clk_period;
		Addr <=  "0010110101010";
		Trees_din <= x"0f005e08";
		wait for Clk_period;
		Addr <=  "0010110101011";
		Trees_din <= x"07ffb104";
		wait for Clk_period;
		Addr <=  "0010110101100";
		Trees_din <= x"ff0417b9";
		wait for Clk_period;
		Addr <=  "0010110101101";
		Trees_din <= x"ffe417b9";
		wait for Clk_period;
		Addr <=  "0010110101110";
		Trees_din <= x"03fce004";
		wait for Clk_period;
		Addr <=  "0010110101111";
		Trees_din <= x"000b17b9";
		wait for Clk_period;
		Addr <=  "0010110110000";
		Trees_din <= x"ff9517b9";
		wait for Clk_period;
		Addr <=  "0010110110001";
		Trees_din <= x"03fdac10";
		wait for Clk_period;
		Addr <=  "0010110110010";
		Trees_din <= x"11014608";
		wait for Clk_period;
		Addr <=  "0010110110011";
		Trees_din <= x"06076c04";
		wait for Clk_period;
		Addr <=  "0010110110100";
		Trees_din <= x"ffe517b9";
		wait for Clk_period;
		Addr <=  "0010110110101";
		Trees_din <= x"006517b9";
		wait for Clk_period;
		Addr <=  "0010110110110";
		Trees_din <= x"1f010e04";
		wait for Clk_period;
		Addr <=  "0010110110111";
		Trees_din <= x"ffd417b9";
		wait for Clk_period;
		Addr <=  "0010110111000";
		Trees_din <= x"011b17b9";
		wait for Clk_period;
		Addr <=  "0010110111001";
		Trees_din <= x"09004708";
		wait for Clk_period;
		Addr <=  "0010110111010";
		Trees_din <= x"01fd6d04";
		wait for Clk_period;
		Addr <=  "0010110111011";
		Trees_din <= x"ffd517b9";
		wait for Clk_period;
		Addr <=  "0010110111100";
		Trees_din <= x"001617b9";
		wait for Clk_period;
		Addr <=  "0010110111101";
		Trees_din <= x"06096c04";
		wait for Clk_period;
		Addr <=  "0010110111110";
		Trees_din <= x"001617b9";
		wait for Clk_period;
		Addr <=  "0010110111111";
		Trees_din <= x"00b517b9";
		wait for Clk_period;
		Addr <=  "0010111000000";
		Trees_din <= x"02fa721c";
		wait for Clk_period;
		Addr <=  "0010111000001";
		Trees_din <= x"01fe3410";
		wait for Clk_period;
		Addr <=  "0010111000010";
		Trees_din <= x"12003f08";
		wait for Clk_period;
		Addr <=  "0010111000011";
		Trees_din <= x"0c010704";
		wait for Clk_period;
		Addr <=  "0010111000100";
		Trees_din <= x"fff717b9";
		wait for Clk_period;
		Addr <=  "0010111000101";
		Trees_din <= x"00d217b9";
		wait for Clk_period;
		Addr <=  "0010111000110";
		Trees_din <= x"0404f704";
		wait for Clk_period;
		Addr <=  "0010111000111";
		Trees_din <= x"003b17b9";
		wait for Clk_period;
		Addr <=  "0010111001000";
		Trees_din <= x"ff9017b9";
		wait for Clk_period;
		Addr <=  "0010111001001";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "0010111001010";
		Trees_din <= x"ff9317b9";
		wait for Clk_period;
		Addr <=  "0010111001011";
		Trees_din <= x"03fe9b04";
		wait for Clk_period;
		Addr <=  "0010111001100";
		Trees_din <= x"00d117b9";
		wait for Clk_period;
		Addr <=  "0010111001101";
		Trees_din <= x"002417b9";
		wait for Clk_period;
		Addr <=  "0010111001110";
		Trees_din <= x"1e023810";
		wait for Clk_period;
		Addr <=  "0010111001111";
		Trees_din <= x"16028108";
		wait for Clk_period;
		Addr <=  "0010111010000";
		Trees_din <= x"1ffec304";
		wait for Clk_period;
		Addr <=  "0010111010001";
		Trees_din <= x"ff8b17b9";
		wait for Clk_period;
		Addr <=  "0010111010010";
		Trees_din <= x"004c17b9";
		wait for Clk_period;
		Addr <=  "0010111010011";
		Trees_din <= x"0b00fe04";
		wait for Clk_period;
		Addr <=  "0010111010100";
		Trees_din <= x"00b917b9";
		wait for Clk_period;
		Addr <=  "0010111010101";
		Trees_din <= x"fff417b9";
		wait for Clk_period;
		Addr <=  "0010111010110";
		Trees_din <= x"06072d08";
		wait for Clk_period;
		Addr <=  "0010111010111";
		Trees_din <= x"12005304";
		wait for Clk_period;
		Addr <=  "0010111011000";
		Trees_din <= x"ff8417b9";
		wait for Clk_period;
		Addr <=  "0010111011001";
		Trees_din <= x"005717b9";
		wait for Clk_period;
		Addr <=  "0010111011010";
		Trees_din <= x"05fe4704";
		wait for Clk_period;
		Addr <=  "0010111011011";
		Trees_din <= x"ff6c17b9";
		wait for Clk_period;
		Addr <=  "0010111011100";
		Trees_din <= x"fff617b9";
		wait for Clk_period;
		Addr <=  "0010111011101";
		Trees_din <= x"03028a04";
		wait for Clk_period;
		Addr <=  "0010111011110";
		Trees_din <= x"008917b9";
		wait for Clk_period;
		Addr <=  "0010111011111";
		Trees_din <= x"060e9010";
		wait for Clk_period;
		Addr <=  "0010111100000";
		Trees_din <= x"08004104";
		wait for Clk_period;
		Addr <=  "0010111100001";
		Trees_din <= x"004317b9";
		wait for Clk_period;
		Addr <=  "0010111100010";
		Trees_din <= x"060dfb04";
		wait for Clk_period;
		Addr <=  "0010111100011";
		Trees_din <= x"002b17b9";
		wait for Clk_period;
		Addr <=  "0010111100100";
		Trees_din <= x"14003b04";
		wait for Clk_period;
		Addr <=  "0010111100101";
		Trees_din <= x"ffed17b9";
		wait for Clk_period;
		Addr <=  "0010111100110";
		Trees_din <= x"ff8a17b9";
		wait for Clk_period;
		Addr <=  "0010111100111";
		Trees_din <= x"0900450c";
		wait for Clk_period;
		Addr <=  "0010111101000";
		Trees_din <= x"04f93c08";
		wait for Clk_period;
		Addr <=  "0010111101001";
		Trees_din <= x"14003b04";
		wait for Clk_period;
		Addr <=  "0010111101010";
		Trees_din <= x"004817b9";
		wait for Clk_period;
		Addr <=  "0010111101011";
		Trees_din <= x"ffff17b9";
		wait for Clk_period;
		Addr <=  "0010111101100";
		Trees_din <= x"007a17b9";
		wait for Clk_period;
		Addr <=  "0010111101101";
		Trees_din <= x"fffe17b9";
		wait for Clk_period;
		Addr <=  "0010111101110";
		Trees_din <= x"0c00e06c";
		wait for Clk_period;
		Addr <=  "0010111101111";
		Trees_din <= x"0d006d34";
		wait for Clk_period;
		Addr <=  "0010111110000";
		Trees_din <= x"1200491c";
		wait for Clk_period;
		Addr <=  "0010111110001";
		Trees_din <= x"09003e0c";
		wait for Clk_period;
		Addr <=  "0010111110010";
		Trees_din <= x"11000004";
		wait for Clk_period;
		Addr <=  "0010111110011";
		Trees_din <= x"ffda195d";
		wait for Clk_period;
		Addr <=  "0010111110100";
		Trees_din <= x"0d006304";
		wait for Clk_period;
		Addr <=  "0010111110101";
		Trees_din <= x"ffdc195d";
		wait for Clk_period;
		Addr <=  "0010111110110";
		Trees_din <= x"00f1195d";
		wait for Clk_period;
		Addr <=  "0010111110111";
		Trees_din <= x"09004208";
		wait for Clk_period;
		Addr <=  "0010111111000";
		Trees_din <= x"15f71604";
		wait for Clk_period;
		Addr <=  "0010111111001";
		Trees_din <= x"0046195d";
		wait for Clk_period;
		Addr <=  "0010111111010";
		Trees_din <= x"ff86195d";
		wait for Clk_period;
		Addr <=  "0010111111011";
		Trees_din <= x"19000104";
		wait for Clk_period;
		Addr <=  "0010111111100";
		Trees_din <= x"00ba195d";
		wait for Clk_period;
		Addr <=  "0010111111101";
		Trees_din <= x"ffb4195d";
		wait for Clk_period;
		Addr <=  "0010111111110";
		Trees_din <= x"12004a0c";
		wait for Clk_period;
		Addr <=  "0010111111111";
		Trees_din <= x"09004208";
		wait for Clk_period;
		Addr <=  "0011000000000";
		Trees_din <= x"13007804";
		wait for Clk_period;
		Addr <=  "0011000000001";
		Trees_din <= x"ffc2195d";
		wait for Clk_period;
		Addr <=  "0011000000010";
		Trees_din <= x"fefa195d";
		wait for Clk_period;
		Addr <=  "0011000000011";
		Trees_din <= x"0079195d";
		wait for Clk_period;
		Addr <=  "0011000000100";
		Trees_din <= x"0407ad08";
		wait for Clk_period;
		Addr <=  "0011000000101";
		Trees_din <= x"08004504";
		wait for Clk_period;
		Addr <=  "0011000000110";
		Trees_din <= x"0050195d";
		wait for Clk_period;
		Addr <=  "0011000000111";
		Trees_din <= x"0006195d";
		wait for Clk_period;
		Addr <=  "0011000001000";
		Trees_din <= x"ff6c195d";
		wait for Clk_period;
		Addr <=  "0011000001001";
		Trees_din <= x"08003d18";
		wait for Clk_period;
		Addr <=  "0011000001010";
		Trees_din <= x"1703ea08";
		wait for Clk_period;
		Addr <=  "0011000001011";
		Trees_din <= x"11005f04";
		wait for Clk_period;
		Addr <=  "0011000001100";
		Trees_din <= x"007c195d";
		wait for Clk_period;
		Addr <=  "0011000001101";
		Trees_din <= x"000a195d";
		wait for Clk_period;
		Addr <=  "0011000001110";
		Trees_din <= x"0a000608";
		wait for Clk_period;
		Addr <=  "0011000001111";
		Trees_din <= x"14003104";
		wait for Clk_period;
		Addr <=  "0011000010000";
		Trees_din <= x"ffba195d";
		wait for Clk_period;
		Addr <=  "0011000010001";
		Trees_din <= x"0060195d";
		wait for Clk_period;
		Addr <=  "0011000010010";
		Trees_din <= x"05fece04";
		wait for Clk_period;
		Addr <=  "0011000010011";
		Trees_din <= x"ff29195d";
		wait for Clk_period;
		Addr <=  "0011000010100";
		Trees_din <= x"ffe3195d";
		wait for Clk_period;
		Addr <=  "0011000010101";
		Trees_din <= x"10000510";
		wait for Clk_period;
		Addr <=  "0011000010110";
		Trees_din <= x"02fa9b08";
		wait for Clk_period;
		Addr <=  "0011000010111";
		Trees_din <= x"01fd4404";
		wait for Clk_period;
		Addr <=  "0011000011000";
		Trees_din <= x"ff96195d";
		wait for Clk_period;
		Addr <=  "0011000011001";
		Trees_din <= x"007d195d";
		wait for Clk_period;
		Addr <=  "0011000011010";
		Trees_din <= x"03015404";
		wait for Clk_period;
		Addr <=  "0011000011011";
		Trees_din <= x"ff8a195d";
		wait for Clk_period;
		Addr <=  "0011000011100";
		Trees_din <= x"0019195d";
		wait for Clk_period;
		Addr <=  "0011000011101";
		Trees_din <= x"1b024608";
		wait for Clk_period;
		Addr <=  "0011000011110";
		Trees_din <= x"0609be04";
		wait for Clk_period;
		Addr <=  "0011000011111";
		Trees_din <= x"ff72195d";
		wait for Clk_period;
		Addr <=  "0011000100000";
		Trees_din <= x"004f195d";
		wait for Clk_period;
		Addr <=  "0011000100001";
		Trees_din <= x"1700c404";
		wait for Clk_period;
		Addr <=  "0011000100010";
		Trees_din <= x"ff68195d";
		wait for Clk_period;
		Addr <=  "0011000100011";
		Trees_din <= x"0027195d";
		wait for Clk_period;
		Addr <=  "0011000100100";
		Trees_din <= x"0c012f38";
		wait for Clk_period;
		Addr <=  "0011000100101";
		Trees_din <= x"07fe5118";
		wait for Clk_period;
		Addr <=  "0011000100110";
		Trees_din <= x"08004e10";
		wait for Clk_period;
		Addr <=  "0011000100111";
		Trees_din <= x"02fd8108";
		wait for Clk_period;
		Addr <=  "0011000101000";
		Trees_din <= x"08004104";
		wait for Clk_period;
		Addr <=  "0011000101001";
		Trees_din <= x"fffe195d";
		wait for Clk_period;
		Addr <=  "0011000101010";
		Trees_din <= x"00a5195d";
		wait for Clk_period;
		Addr <=  "0011000101011";
		Trees_din <= x"08004a04";
		wait for Clk_period;
		Addr <=  "0011000101100";
		Trees_din <= x"ff99195d";
		wait for Clk_period;
		Addr <=  "0011000101101";
		Trees_din <= x"0069195d";
		wait for Clk_period;
		Addr <=  "0011000101110";
		Trees_din <= x"1b027004";
		wait for Clk_period;
		Addr <=  "0011000101111";
		Trees_din <= x"ff1c195d";
		wait for Clk_period;
		Addr <=  "0011000110000";
		Trees_din <= x"001f195d";
		wait for Clk_period;
		Addr <=  "0011000110001";
		Trees_din <= x"04054b10";
		wait for Clk_period;
		Addr <=  "0011000110010";
		Trees_din <= x"11000208";
		wait for Clk_period;
		Addr <=  "0011000110011";
		Trees_din <= x"0c012704";
		wait for Clk_period;
		Addr <=  "0011000110100";
		Trees_din <= x"0082195d";
		wait for Clk_period;
		Addr <=  "0011000110101";
		Trees_din <= x"ff81195d";
		wait for Clk_period;
		Addr <=  "0011000110110";
		Trees_din <= x"11000604";
		wait for Clk_period;
		Addr <=  "0011000110111";
		Trees_din <= x"fed7195d";
		wait for Clk_period;
		Addr <=  "0011000111000";
		Trees_din <= x"ffa3195d";
		wait for Clk_period;
		Addr <=  "0011000111001";
		Trees_din <= x"05fe3508";
		wait for Clk_period;
		Addr <=  "0011000111010";
		Trees_din <= x"1b025104";
		wait for Clk_period;
		Addr <=  "0011000111011";
		Trees_din <= x"ff38195d";
		wait for Clk_period;
		Addr <=  "0011000111100";
		Trees_din <= x"fffa195d";
		wait for Clk_period;
		Addr <=  "0011000111101";
		Trees_din <= x"06082604";
		wait for Clk_period;
		Addr <=  "0011000111110";
		Trees_din <= x"0021195d";
		wait for Clk_period;
		Addr <=  "0011000111111";
		Trees_din <= x"00c8195d";
		wait for Clk_period;
		Addr <=  "0011001000000";
		Trees_din <= x"15f71a10";
		wait for Clk_period;
		Addr <=  "0011001000001";
		Trees_din <= x"11000008";
		wait for Clk_period;
		Addr <=  "0011001000010";
		Trees_din <= x"0f005604";
		wait for Clk_period;
		Addr <=  "0011001000011";
		Trees_din <= x"ffcd195d";
		wait for Clk_period;
		Addr <=  "0011001000100";
		Trees_din <= x"00c7195d";
		wait for Clk_period;
		Addr <=  "0011001000101";
		Trees_din <= x"08004c04";
		wait for Clk_period;
		Addr <=  "0011001000110";
		Trees_din <= x"ff09195d";
		wait for Clk_period;
		Addr <=  "0011001000111";
		Trees_din <= x"ffc7195d";
		wait for Clk_period;
		Addr <=  "0011001001000";
		Trees_din <= x"0c013710";
		wait for Clk_period;
		Addr <=  "0011001001001";
		Trees_din <= x"1afcd008";
		wait for Clk_period;
		Addr <=  "0011001001010";
		Trees_din <= x"11000804";
		wait for Clk_period;
		Addr <=  "0011001001011";
		Trees_din <= x"0030195d";
		wait for Clk_period;
		Addr <=  "0011001001100";
		Trees_din <= x"00ee195d";
		wait for Clk_period;
		Addr <=  "0011001001101";
		Trees_din <= x"11001004";
		wait for Clk_period;
		Addr <=  "0011001001110";
		Trees_din <= x"0072195d";
		wait for Clk_period;
		Addr <=  "0011001001111";
		Trees_din <= x"ff28195d";
		wait for Clk_period;
		Addr <=  "0011001010000";
		Trees_din <= x"10008a08";
		wait for Clk_period;
		Addr <=  "0011001010001";
		Trees_din <= x"01fd3604";
		wait for Clk_period;
		Addr <=  "0011001010010";
		Trees_din <= x"ffe5195d";
		wait for Clk_period;
		Addr <=  "0011001010011";
		Trees_din <= x"0042195d";
		wait for Clk_period;
		Addr <=  "0011001010100";
		Trees_din <= x"1000d004";
		wait for Clk_period;
		Addr <=  "0011001010101";
		Trees_din <= x"ffc2195d";
		wait for Clk_period;
		Addr <=  "0011001010110";
		Trees_din <= x"000a195d";
		wait for Clk_period;
		Addr <=  "0011001010111";
		Trees_din <= x"00026268";
		wait for Clk_period;
		Addr <=  "0011001011000";
		Trees_din <= x"060c1740";
		wait for Clk_period;
		Addr <=  "0011001011001";
		Trees_din <= x"1703e520";
		wait for Clk_period;
		Addr <=  "0011001011010";
		Trees_din <= x"1703d010";
		wait for Clk_period;
		Addr <=  "0011001011011";
		Trees_din <= x"060be908";
		wait for Clk_period;
		Addr <=  "0011001011100";
		Trees_din <= x"12004604";
		wait for Clk_period;
		Addr <=  "0011001011101";
		Trees_din <= x"00121a31";
		wait for Clk_period;
		Addr <=  "0011001011110";
		Trees_din <= x"fff11a31";
		wait for Clk_period;
		Addr <=  "0011001011111";
		Trees_din <= x"05fe6e04";
		wait for Clk_period;
		Addr <=  "0011001100000";
		Trees_din <= x"00321a31";
		wait for Clk_period;
		Addr <=  "0011001100001";
		Trees_din <= x"fef01a31";
		wait for Clk_period;
		Addr <=  "0011001100010";
		Trees_din <= x"00fd4808";
		wait for Clk_period;
		Addr <=  "0011001100011";
		Trees_din <= x"060af404";
		wait for Clk_period;
		Addr <=  "0011001100100";
		Trees_din <= x"ff501a31";
		wait for Clk_period;
		Addr <=  "0011001100101";
		Trees_din <= x"00641a31";
		wait for Clk_period;
		Addr <=  "0011001100110";
		Trees_din <= x"0d008904";
		wait for Clk_period;
		Addr <=  "0011001100111";
		Trees_din <= x"00031a31";
		wait for Clk_period;
		Addr <=  "0011001101000";
		Trees_din <= x"ff7f1a31";
		wait for Clk_period;
		Addr <=  "0011001101001";
		Trees_din <= x"1703ec10";
		wait for Clk_period;
		Addr <=  "0011001101010";
		Trees_din <= x"0e002a08";
		wait for Clk_period;
		Addr <=  "0011001101011";
		Trees_din <= x"03014204";
		wait for Clk_period;
		Addr <=  "0011001101100";
		Trees_din <= x"00b51a31";
		wait for Clk_period;
		Addr <=  "0011001101101";
		Trees_din <= x"ffb41a31";
		wait for Clk_period;
		Addr <=  "0011001101110";
		Trees_din <= x"02fa5504";
		wait for Clk_period;
		Addr <=  "0011001101111";
		Trees_din <= x"ff651a31";
		wait for Clk_period;
		Addr <=  "0011001110000";
		Trees_din <= x"004e1a31";
		wait for Clk_period;
		Addr <=  "0011001110001";
		Trees_din <= x"10013308";
		wait for Clk_period;
		Addr <=  "0011001110010";
		Trees_din <= x"01feff04";
		wait for Clk_period;
		Addr <=  "0011001110011";
		Trees_din <= x"00041a31";
		wait for Clk_period;
		Addr <=  "0011001110100";
		Trees_din <= x"00621a31";
		wait for Clk_period;
		Addr <=  "0011001110101";
		Trees_din <= x"060a4e04";
		wait for Clk_period;
		Addr <=  "0011001110110";
		Trees_din <= x"ff5e1a31";
		wait for Clk_period;
		Addr <=  "0011001110111";
		Trees_din <= x"00231a31";
		wait for Clk_period;
		Addr <=  "0011001111000";
		Trees_din <= x"10000210";
		wait for Clk_period;
		Addr <=  "0011001111001";
		Trees_din <= x"08004304";
		wait for Clk_period;
		Addr <=  "0011001111010";
		Trees_din <= x"ff201a31";
		wait for Clk_period;
		Addr <=  "0011001111011";
		Trees_din <= x"08005108";
		wait for Clk_period;
		Addr <=  "0011001111100";
		Trees_din <= x"00fec404";
		wait for Clk_period;
		Addr <=  "0011001111101";
		Trees_din <= x"00691a31";
		wait for Clk_period;
		Addr <=  "0011001111110";
		Trees_din <= x"000d1a31";
		wait for Clk_period;
		Addr <=  "0011001111111";
		Trees_din <= x"ff7a1a31";
		wait for Clk_period;
		Addr <=  "0011010000000";
		Trees_din <= x"07feb710";
		wait for Clk_period;
		Addr <=  "0011010000001";
		Trees_din <= x"1c026208";
		wait for Clk_period;
		Addr <=  "0011010000010";
		Trees_din <= x"0b010104";
		wait for Clk_period;
		Addr <=  "0011010000011";
		Trees_din <= x"00891a31";
		wait for Clk_period;
		Addr <=  "0011010000100";
		Trees_din <= x"ff7d1a31";
		wait for Clk_period;
		Addr <=  "0011010000101";
		Trees_din <= x"08004504";
		wait for Clk_period;
		Addr <=  "0011010000110";
		Trees_din <= x"002f1a31";
		wait for Clk_period;
		Addr <=  "0011010000111";
		Trees_din <= x"ffc81a31";
		wait for Clk_period;
		Addr <=  "0011010001000";
		Trees_din <= x"07014504";
		wait for Clk_period;
		Addr <=  "0011010001001";
		Trees_din <= x"00941a31";
		wait for Clk_period;
		Addr <=  "0011010001010";
		Trees_din <= x"001c1a31";
		wait for Clk_period;
		Addr <=  "0011010001011";
		Trees_din <= x"ff881a31";
		wait for Clk_period;
		Addr <=  "0011010001100";
		Trees_din <= x"06013010";
		wait for Clk_period;
		Addr <=  "0011010001101";
		Trees_din <= x"1300ce08";
		wait for Clk_period;
		Addr <=  "0011010001110";
		Trees_din <= x"09004d04";
		wait for Clk_period;
		Addr <=  "0011010001111";
		Trees_din <= x"ff771b3d";
		wait for Clk_period;
		Addr <=  "0011010010000";
		Trees_din <= x"00261b3d";
		wait for Clk_period;
		Addr <=  "0011010010001";
		Trees_din <= x"0f008504";
		wait for Clk_period;
		Addr <=  "0011010010010";
		Trees_din <= x"00651b3d";
		wait for Clk_period;
		Addr <=  "0011010010011";
		Trees_din <= x"ffaf1b3d";
		wait for Clk_period;
		Addr <=  "0011010010100";
		Trees_din <= x"05fcb938";
		wait for Clk_period;
		Addr <=  "0011010010101";
		Trees_din <= x"02fa7c1c";
		wait for Clk_period;
		Addr <=  "0011010010110";
		Trees_din <= x"05fc2c10";
		wait for Clk_period;
		Addr <=  "0011010010111";
		Trees_din <= x"18005a08";
		wait for Clk_period;
		Addr <=  "0011010011000";
		Trees_din <= x"1300c604";
		wait for Clk_period;
		Addr <=  "0011010011001";
		Trees_din <= x"ffd51b3d";
		wait for Clk_period;
		Addr <=  "0011010011010";
		Trees_din <= x"00761b3d";
		wait for Clk_period;
		Addr <=  "0011010011011";
		Trees_din <= x"03fa3e04";
		wait for Clk_period;
		Addr <=  "0011010011100";
		Trees_din <= x"00071b3d";
		wait for Clk_period;
		Addr <=  "0011010011101";
		Trees_din <= x"ff4a1b3d";
		wait for Clk_period;
		Addr <=  "0011010011110";
		Trees_din <= x"0f006504";
		wait for Clk_period;
		Addr <=  "0011010011111";
		Trees_din <= x"00b91b3d";
		wait for Clk_period;
		Addr <=  "0011010100000";
		Trees_din <= x"07007a04";
		wait for Clk_period;
		Addr <=  "0011010100001";
		Trees_din <= x"ff8b1b3d";
		wait for Clk_period;
		Addr <=  "0011010100010";
		Trees_din <= x"00261b3d";
		wait for Clk_period;
		Addr <=  "0011010100011";
		Trees_din <= x"0d00670c";
		wait for Clk_period;
		Addr <=  "0011010100100";
		Trees_din <= x"0c02c508";
		wait for Clk_period;
		Addr <=  "0011010100101";
		Trees_din <= x"01fd9004";
		wait for Clk_period;
		Addr <=  "0011010100110";
		Trees_din <= x"ff611b3d";
		wait for Clk_period;
		Addr <=  "0011010100111";
		Trees_din <= x"00151b3d";
		wait for Clk_period;
		Addr <=  "0011010101000";
		Trees_din <= x"00c31b3d";
		wait for Clk_period;
		Addr <=  "0011010101001";
		Trees_din <= x"12003d08";
		wait for Clk_period;
		Addr <=  "0011010101010";
		Trees_din <= x"18004e04";
		wait for Clk_period;
		Addr <=  "0011010101011";
		Trees_din <= x"00661b3d";
		wait for Clk_period;
		Addr <=  "0011010101100";
		Trees_din <= x"ff8e1b3d";
		wait for Clk_period;
		Addr <=  "0011010101101";
		Trees_din <= x"1300ab04";
		wait for Clk_period;
		Addr <=  "0011010101110";
		Trees_din <= x"002e1b3d";
		wait for Clk_period;
		Addr <=  "0011010101111";
		Trees_din <= x"00a51b3d";
		wait for Clk_period;
		Addr <=  "0011010110000";
		Trees_din <= x"02fa7c20";
		wait for Clk_period;
		Addr <=  "0011010110001";
		Trees_din <= x"09004010";
		wait for Clk_period;
		Addr <=  "0011010110010";
		Trees_din <= x"00fcdd08";
		wait for Clk_period;
		Addr <=  "0011010110011";
		Trees_din <= x"01fd5c04";
		wait for Clk_period;
		Addr <=  "0011010110100";
		Trees_din <= x"ff591b3d";
		wait for Clk_period;
		Addr <=  "0011010110101";
		Trees_din <= x"00121b3d";
		wait for Clk_period;
		Addr <=  "0011010110110";
		Trees_din <= x"12003304";
		wait for Clk_period;
		Addr <=  "0011010110111";
		Trees_din <= x"ffb11b3d";
		wait for Clk_period;
		Addr <=  "0011010111000";
		Trees_din <= x"005c1b3d";
		wait for Clk_period;
		Addr <=  "0011010111001";
		Trees_din <= x"1afc4f08";
		wait for Clk_period;
		Addr <=  "0011010111010";
		Trees_din <= x"0f008104";
		wait for Clk_period;
		Addr <=  "0011010111011";
		Trees_din <= x"ff9f1b3d";
		wait for Clk_period;
		Addr <=  "0011010111100";
		Trees_din <= x"002a1b3d";
		wait for Clk_period;
		Addr <=  "0011010111101";
		Trees_din <= x"1703dc04";
		wait for Clk_period;
		Addr <=  "0011010111110";
		Trees_din <= x"009a1b3d";
		wait for Clk_period;
		Addr <=  "0011010111111";
		Trees_din <= x"ffce1b3d";
		wait for Clk_period;
		Addr <=  "0011011000000";
		Trees_din <= x"0d005f10";
		wait for Clk_period;
		Addr <=  "0011011000001";
		Trees_din <= x"07010608";
		wait for Clk_period;
		Addr <=  "0011011000010";
		Trees_din <= x"0f005d04";
		wait for Clk_period;
		Addr <=  "0011011000011";
		Trees_din <= x"ffda1b3d";
		wait for Clk_period;
		Addr <=  "0011011000100";
		Trees_din <= x"00541b3d";
		wait for Clk_period;
		Addr <=  "0011011000101";
		Trees_din <= x"03fb7b04";
		wait for Clk_period;
		Addr <=  "0011011000110";
		Trees_din <= x"ffcf1b3d";
		wait for Clk_period;
		Addr <=  "0011011000111";
		Trees_din <= x"00d81b3d";
		wait for Clk_period;
		Addr <=  "0011011001000";
		Trees_din <= x"13010908";
		wait for Clk_period;
		Addr <=  "0011011001001";
		Trees_din <= x"0401c404";
		wait for Clk_period;
		Addr <=  "0011011001010";
		Trees_din <= x"000e1b3d";
		wait for Clk_period;
		Addr <=  "0011011001011";
		Trees_din <= x"ffe71b3d";
		wait for Clk_period;
		Addr <=  "0011011001100";
		Trees_din <= x"05ff2204";
		wait for Clk_period;
		Addr <=  "0011011001101";
		Trees_din <= x"00921b3d";
		wait for Clk_period;
		Addr <=  "0011011001110";
		Trees_din <= x"fff41b3d";
		wait for Clk_period;
		Addr <=  "0011011001111";
		Trees_din <= x"0605f45c";
		wait for Clk_period;
		Addr <=  "0011011010000";
		Trees_din <= x"0f007e3c";
		wait for Clk_period;
		Addr <=  "0011011010001";
		Trees_din <= x"0f007420";
		wait for Clk_period;
		Addr <=  "0011011010010";
		Trees_din <= x"18007810";
		wait for Clk_period;
		Addr <=  "0011011010011";
		Trees_din <= x"08004308";
		wait for Clk_period;
		Addr <=  "0011011010100";
		Trees_din <= x"17033804";
		wait for Clk_period;
		Addr <=  "0011011010101";
		Trees_din <= x"ffb91c91";
		wait for Clk_period;
		Addr <=  "0011011010110";
		Trees_din <= x"009f1c91";
		wait for Clk_period;
		Addr <=  "0011011010111";
		Trees_din <= x"01fe3204";
		wait for Clk_period;
		Addr <=  "0011011011000";
		Trees_din <= x"ff781c91";
		wait for Clk_period;
		Addr <=  "0011011011001";
		Trees_din <= x"000e1c91";
		wait for Clk_period;
		Addr <=  "0011011011010";
		Trees_din <= x"0e005208";
		wait for Clk_period;
		Addr <=  "0011011011011";
		Trees_din <= x"09004904";
		wait for Clk_period;
		Addr <=  "0011011011100";
		Trees_din <= x"ff971c91";
		wait for Clk_period;
		Addr <=  "0011011011101";
		Trees_din <= x"007d1c91";
		wait for Clk_period;
		Addr <=  "0011011011110";
		Trees_din <= x"03026804";
		wait for Clk_period;
		Addr <=  "0011011011111";
		Trees_din <= x"fff31c91";
		wait for Clk_period;
		Addr <=  "0011011100000";
		Trees_din <= x"009f1c91";
		wait for Clk_period;
		Addr <=  "0011011100001";
		Trees_din <= x"00fd980c";
		wait for Clk_period;
		Addr <=  "0011011100010";
		Trees_din <= x"05fd3a08";
		wait for Clk_period;
		Addr <=  "0011011100011";
		Trees_din <= x"03fc2604";
		wait for Clk_period;
		Addr <=  "0011011100100";
		Trees_din <= x"ffe11c91";
		wait for Clk_period;
		Addr <=  "0011011100101";
		Trees_din <= x"01021c91";
		wait for Clk_period;
		Addr <=  "0011011100110";
		Trees_din <= x"ff811c91";
		wait for Clk_period;
		Addr <=  "0011011100111";
		Trees_din <= x"18008508";
		wait for Clk_period;
		Addr <=  "0011011101000";
		Trees_din <= x"1602bc04";
		wait for Clk_period;
		Addr <=  "0011011101001";
		Trees_din <= x"00191c91";
		wait for Clk_period;
		Addr <=  "0011011101010";
		Trees_din <= x"ff711c91";
		wait for Clk_period;
		Addr <=  "0011011101011";
		Trees_din <= x"10012f04";
		wait for Clk_period;
		Addr <=  "0011011101100";
		Trees_din <= x"ff9f1c91";
		wait for Clk_period;
		Addr <=  "0011011101101";
		Trees_din <= x"008f1c91";
		wait for Clk_period;
		Addr <=  "0011011101110";
		Trees_din <= x"1300d418";
		wait for Clk_period;
		Addr <=  "0011011101111";
		Trees_din <= x"1000b60c";
		wait for Clk_period;
		Addr <=  "0011011110000";
		Trees_din <= x"1afc5408";
		wait for Clk_period;
		Addr <=  "0011011110001";
		Trees_din <= x"0c009104";
		wait for Clk_period;
		Addr <=  "0011011110010";
		Trees_din <= x"009f1c91";
		wait for Clk_period;
		Addr <=  "0011011110011";
		Trees_din <= x"ffd11c91";
		wait for Clk_period;
		Addr <=  "0011011110100";
		Trees_din <= x"ff6f1c91";
		wait for Clk_period;
		Addr <=  "0011011110101";
		Trees_din <= x"0408ab08";
		wait for Clk_period;
		Addr <=  "0011011110110";
		Trees_din <= x"02fcc604";
		wait for Clk_period;
		Addr <=  "0011011110111";
		Trees_din <= x"00cb1c91";
		wait for Clk_period;
		Addr <=  "0011011111000";
		Trees_din <= x"ffd51c91";
		wait for Clk_period;
		Addr <=  "0011011111001";
		Trees_din <= x"ff981c91";
		wait for Clk_period;
		Addr <=  "0011011111010";
		Trees_din <= x"15f79d04";
		wait for Clk_period;
		Addr <=  "0011011111011";
		Trees_din <= x"00281c91";
		wait for Clk_period;
		Addr <=  "0011011111100";
		Trees_din <= x"ff6f1c91";
		wait for Clk_period;
		Addr <=  "0011011111101";
		Trees_din <= x"03fa2d18";
		wait for Clk_period;
		Addr <=  "0011011111110";
		Trees_din <= x"0b00ba0c";
		wait for Clk_period;
		Addr <=  "0011011111111";
		Trees_din <= x"08004f08";
		wait for Clk_period;
		Addr <=  "0011100000000";
		Trees_din <= x"04050804";
		wait for Clk_period;
		Addr <=  "0011100000001";
		Trees_din <= x"00631c91";
		wait for Clk_period;
		Addr <=  "0011100000010";
		Trees_din <= x"ff351c91";
		wait for Clk_period;
		Addr <=  "0011100000011";
		Trees_din <= x"00cb1c91";
		wait for Clk_period;
		Addr <=  "0011100000100";
		Trees_din <= x"06088308";
		wait for Clk_period;
		Addr <=  "0011100000101";
		Trees_din <= x"10007f04";
		wait for Clk_period;
		Addr <=  "0011100000110";
		Trees_din <= x"00751c91";
		wait for Clk_period;
		Addr <=  "0011100000111";
		Trees_din <= x"ff9d1c91";
		wait for Clk_period;
		Addr <=  "0011100001000";
		Trees_din <= x"00c71c91";
		wait for Clk_period;
		Addr <=  "0011100001001";
		Trees_din <= x"13010920";
		wait for Clk_period;
		Addr <=  "0011100001010";
		Trees_din <= x"0e002310";
		wait for Clk_period;
		Addr <=  "0011100001011";
		Trees_din <= x"02fb0308";
		wait for Clk_period;
		Addr <=  "0011100001100";
		Trees_din <= x"05fdf904";
		wait for Clk_period;
		Addr <=  "0011100001101";
		Trees_din <= x"fff51c91";
		wait for Clk_period;
		Addr <=  "0011100001110";
		Trees_din <= x"006e1c91";
		wait for Clk_period;
		Addr <=  "0011100001111";
		Trees_din <= x"04020c04";
		wait for Clk_period;
		Addr <=  "0011100010000";
		Trees_din <= x"00181c91";
		wait for Clk_period;
		Addr <=  "0011100010001";
		Trees_din <= x"ff9d1c91";
		wait for Clk_period;
		Addr <=  "0011100010010";
		Trees_din <= x"0c000708";
		wait for Clk_period;
		Addr <=  "0011100010011";
		Trees_din <= x"18009804";
		wait for Clk_period;
		Addr <=  "0011100010100";
		Trees_din <= x"006a1c91";
		wait for Clk_period;
		Addr <=  "0011100010101";
		Trees_din <= x"ffe31c91";
		wait for Clk_period;
		Addr <=  "0011100010110";
		Trees_din <= x"10000504";
		wait for Clk_period;
		Addr <=  "0011100010111";
		Trees_din <= x"ffc11c91";
		wait for Clk_period;
		Addr <=  "0011100011000";
		Trees_din <= x"00081c91";
		wait for Clk_period;
		Addr <=  "0011100011001";
		Trees_din <= x"1c026108";
		wait for Clk_period;
		Addr <=  "0011100011010";
		Trees_din <= x"08003c04";
		wait for Clk_period;
		Addr <=  "0011100011011";
		Trees_din <= x"ff801c91";
		wait for Clk_period;
		Addr <=  "0011100011100";
		Trees_din <= x"001a1c91";
		wait for Clk_period;
		Addr <=  "0011100011101";
		Trees_din <= x"060bc308";
		wait for Clk_period;
		Addr <=  "0011100011110";
		Trees_din <= x"05ff0804";
		wait for Clk_period;
		Addr <=  "0011100011111";
		Trees_din <= x"00b01c91";
		wait for Clk_period;
		Addr <=  "0011100100000";
		Trees_din <= x"fffc1c91";
		wait for Clk_period;
		Addr <=  "0011100100001";
		Trees_din <= x"0c016104";
		wait for Clk_period;
		Addr <=  "0011100100010";
		Trees_din <= x"00431c91";
		wait for Clk_period;
		Addr <=  "0011100100011";
		Trees_din <= x"ff951c91";
		wait for Clk_period;
		Addr <=  "0011100100100";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  1
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"0406846c";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"04045e30";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"04016f10";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"1a051c0c";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"12002a04";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"000f016d";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"0d00bd04";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"ff5d016d";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"0000016d";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"0037016d";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"03ffdb10";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"04038108";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"0c031404";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"ff7c016d";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"0031016d";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"1afa3e04";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"0065016d";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"ffbd016d";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"06090c08";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"0603f604";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"ffb2016d";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"0103016d";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"07fe6c04";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"ff84016d";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"007b016d";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"060af420";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"0701d110";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"06082608";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"01ff7704";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"01d0016d";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"ffc7016d";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"07001f04";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"0103016d";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"0020016d";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"07062508";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"04056704";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"ffce016d";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"00a1016d";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"15f73704";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"000f016d";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"ff60016d";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"0f007f0c";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"10000004";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"0089016d";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"08003e04";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"fff0016d";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"ff58016d";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"05fd6f08";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"07fe0304";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"0037016d";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"0235016d";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"12004d04";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"ff87016d";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"012b016d";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"0408c134";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"0705471c";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"01fea90c";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"1a013e08";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"1af8d904";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"0093016d";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"0312016d";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"fff3016d";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"04077208";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"02fb0e04";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"ffc1016d";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"0127016d";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"01006304";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"02d1016d";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"ff88016d";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"1c026b10";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"07072708";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"03fb3804";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"0037016d";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"02e7016d";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"0001c404";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"ffa4016d";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"0037016d";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"05fbb604";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"0089016d";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"ff6d016d";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"07079b0c";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"0607fe08";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"01044c04";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"0435016d";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"014f016d";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"00ca016d";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"040bfb04";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"ff7c016d";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"070a2304";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"0235016d";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"0037016d";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"0405835c";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"0401d21c";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"1a051c18";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"04016f0c";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"12002a04";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"001902c1";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"0d00bd04";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"ff6502c1";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"000e02c1";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"15f70004";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"013b02c1";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"02ff3904";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"ff6902c1";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"007e02c1";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"003c02c1";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"060bc320";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"0701d110";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"0609be08";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"08005204";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"008402c1";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"ff7902c1";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"0404f704";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"ffe402c1";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"007b02c1";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"0d005f08";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"0e004d04";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"00f002c1";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"ff8702c1";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"09004c04";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"ff8102c1";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"007f02c1";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"05fd3a10";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"03fc1008";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"1afb4e04";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"003602c1";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"015f02c1";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"11011404";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"ff7802c1";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"003d02c1";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"10000508";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"14003d04";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"015302c1";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"ff7902c1";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"0f005d04";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"003f02c1";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"ff6202c1";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"04075a34";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"03feef20";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"01feae10";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"00005008";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"ffc602c1";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"010c02c1";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"11000104";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"016c02c1";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"ff9f02c1";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"15fa9408";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"03fe4f04";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"ffd602c1";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"011802c1";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"03fc7804";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"026e02c1";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"000702c1";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"0e002008";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"07006e04";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"ff8502c1";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"00d902c1";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"0f005d04";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"ffa402c1";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"01fff104";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"021902c1";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"003302c1";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"0003ad14";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"040b2b10";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"01ffb308";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"0702cf04";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"019a02c1";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"011a02c1";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"03fd8304";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"003a02c1";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"016b02c1";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"01c702c1";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"0f007004";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"003c02c1";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"ff7102c1";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"04056750";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"0401d218";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"04fb9604";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"ff5b042d";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"03004a04";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"ff5c042d";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"04014a08";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"03008104";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"005d042d";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"ff81042d";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"01fd8404";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"00e4042d";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"ffb7042d";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"060c0f20";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"0701dd10";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"01fd9608";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"03fc7804";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"00c7042d";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"0038042d";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"0d006d04";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"ffbe042d";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"002e042d";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"0d005f08";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"03fdca04";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"00c3042d";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"ff8c042d";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"09004d04";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"ff81042d";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"005e042d";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"08005410";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"08003a08";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"0e003304";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"ff9e042d";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"00db042d";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"0b010604";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"ff5d042d";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"000d042d";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"05fdc604";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"0145042d";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"ff97042d";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"0406cb40";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"07021920";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"060a4110";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"03fae008";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"ffe6042d";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"0190042d";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"1f026f04";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"007f042d";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"0104042d";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"02fb6b08";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"07feb004";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"ffd3042d";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"00de042d";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"0c002104";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"0032042d";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"ff5e042d";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"1c028210";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"01fd6508";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"11001604";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"00e7042d";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"ff79042d";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"03fec304";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"ff71042d";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"0087042d";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"0704b808";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"04068404";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"018c042d";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"ffd9042d";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"09004704";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"ff8f042d";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"003f042d";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"0003ad20";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"06087510";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"07081908";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"040b2b04";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"00fd042d";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"013c042d";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"00028c04";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"ff9e042d";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"0122042d";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"10007608";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"08004504";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"ff9b042d";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"00ad042d";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"00fd4004";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"0002042d";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"0146042d";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"0d006504";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"0036042d";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"ff75042d";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"0404c960";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"04016f2c";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"11028920";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"09004a10";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"19008308";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"0b012704";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"ff670589";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"00190589";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"10006404";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"00dd0589";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"ff840589";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"0c027108";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"01fc5a04";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"00310589";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"ff6c0589";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"1300ae04";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"ffa40589";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"01640589";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"04fe2504";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"ff7e0589";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"04000604";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"01410589";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"ffa90589";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"060ae620";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"0701dd10";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"10036e08";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"1af8d904";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"015e0589";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"00150589";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"08004404";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"00370589";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"02440589";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"0e004908";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"00fed004";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"ffc90589";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"ff5f0589";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"14004c04";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"00d80589";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"ffa30589";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"0c034410";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"08005908";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"0f009d04";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"ff900589";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"00830589";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"03fca004";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"015c0589";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"ff980589";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"00c10589";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"0406cb24";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"0c000710";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"0700a90c";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"0b00fe08";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"0b007404";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"00e60589";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"ff970589";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"012a0589";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"ff5a0589";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"060c2410";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"0703b108";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"01fcdb04";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"00e40589";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"00700589";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"0f008904";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"ffbd0589";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"00b90589";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"ff760589";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"040b2b1c";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"0100bd10";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"07072708";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"10038204";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"00c00589";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"00000589";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"15f7ad04";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"00440589";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"ff720589";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"18005504";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"00a70589";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"19000704";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"ff4c0589";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"002f0589";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"070a230c";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"07fbb604";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"005d0589";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"0b011504";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"00fe0589";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"00690589";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"fffd0589";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"04042e68";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"04016f2c";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"11028920";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"09004a10";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"19008308";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"0b012704";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"ff6c0725";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"00190725";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"07feb004";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"ff8a0725";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"00d60725";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"0c027108";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"11000204";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"00410725";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"ff700725";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"14004704";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"01640725";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"ffa30725";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"04fe2504";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"ff850725";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"1b026104";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"010c0725";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"ffac0725";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"03ffdb1c";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"0c02e210";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"03fcf208";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"0f006904";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"00e10725";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"ffc90725";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"09002404";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"008e0725";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"ff8a0725";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"03fcb204";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"ff750725";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"19000104";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"ffcf0725";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"013e0725";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"01fe3410";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"0a000e08";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"0e002c04";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"00590725";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"ff6d0725";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"03016c04";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"01010725";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"00130725";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"08004608";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"1602fc04";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"002b0725";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"ff5f0725";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"18007404";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"00f80725";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"ff830725";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"04068428";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"09004c14";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"12005c10";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"00001f08";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"01fc7404";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"00e90725";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"00430725";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"0c013c04";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"003b0725";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"ff580725";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"ff5f0725";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"1f02830c";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"08005408";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"19000a04";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"01ea0725";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"00100725";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"ff9e0725";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"16018204";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"00340725";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"ff7e0725";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"04095320";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"03fdb210";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"01ffb308";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"0702cf04";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"008c0725";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"003c0725";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"19001c04";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"ff930725";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"00fc0725";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"1b028708";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"09003104";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"ffb40725";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"00e40725";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"00fedc04";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"ff560725";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"fff50725";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"0705d210";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"05fd2e08";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"10036e04";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"00db0725";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"000e0725";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"0b006504";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"ffd90725";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"00ad0725";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"040b0008";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"0a00e304";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"ff450725";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"00350725";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"0a027904";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"00cf0725";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"ff9c0725";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"04042e50";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"04016f20";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"1af8eb08";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"0c018504";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"00d70871";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"ff9d0871";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"1ffd6208";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"0b00e804";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"ff960871";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"00bc0871";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"09004a08";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"0f006504";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"ffc30871";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"ff6e0871";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"0c027104";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"ff950871";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"009a0871";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"03ffdb1c";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"0c02e210";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"03fcf208";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"07ff8904";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"006c0871";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"ffb80871";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"09002404";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"007d0871";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"ff930871";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"03fcb204";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"ff7c0871";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"0d007e04";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"00e30871";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"ff980871";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"1af8c104";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"01770871";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"03030708";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"0d006604";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"ffa70871";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"00700871";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"11000004";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"00820871";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"ff790871";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"0408c120";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"00031a1c";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"060b2c10";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"07001f08";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"01fedd04";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"00800871";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"00200871";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"06082604";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"004f0871";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"fffa0871";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"03fcb208";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"0f007f04";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"ffe30871";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"00d40871";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"ff640871";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"ff6e0871";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"08005020";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"17040010";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"070a2308";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"0e002704";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"00880871";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"00c10871";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"0b00b304";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"ffa40871";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"00340871";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"05fcca08";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"08004a04";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"00c80871";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"00210871";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"01feb604";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"00810871";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"ff580871";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"0d008a10";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"040b2b08";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"01fe2e04";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"00160871";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"ff080871";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"0703b104";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"00bf0871";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"ffe70871";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"12006604";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"00cd0871";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"002c0871";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"0404b548";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"04016f20";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"04fb9604";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"ff6509e1";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"01feb60c";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"05053c08";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"1af8eb04";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"008509e1";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"ff7b09e1";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"00be09e1";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"01fef208";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"18006604";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"ffad09e1";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"016309e1";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"09004a04";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"ff7509e1";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"00a609e1";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"01fb8f08";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"0402d004";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"001d09e1";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"019e09e1";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"07020e10";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"060c0f08";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"0a000304";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"009b09e1";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"000709e1";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"05fd2a04";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"009c09e1";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"ff8609e1";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"0d006308";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"0b00c104";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"010009e1";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"ff8009e1";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"16040004";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"ff6309e1";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"ffb809e1";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"04095338";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"07004720";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"05fd8d10";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"00feb608";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"03fc3404";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"00c609e1";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"005409e1";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"06085504";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"008009e1";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"ffc809e1";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"08003d08";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"00fd8204";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"014509e1";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"005109e1";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"05fdba04";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"ffc709e1";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"003e09e1";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"0f009d10";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"04066f08";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"05fd0504";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"ffc309e1";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"002f09e1";
		wait for Clk_period;
		Addr <=  "0001001010111";
		Trees_din <= x"10001104";
		wait for Clk_period;
		Addr <=  "0001001011000";
		Trees_din <= x"00b009e1";
		wait for Clk_period;
		Addr <=  "0001001011001";
		Trees_din <= x"003209e1";
		wait for Clk_period;
		Addr <=  "0001001011010";
		Trees_din <= x"06005804";
		wait for Clk_period;
		Addr <=  "0001001011011";
		Trees_din <= x"005809e1";
		wait for Clk_period;
		Addr <=  "0001001011100";
		Trees_din <= x"012d09e1";
		wait for Clk_period;
		Addr <=  "0001001011101";
		Trees_din <= x"07041c1c";
		wait for Clk_period;
		Addr <=  "0001001011110";
		Trees_din <= x"0f00660c";
		wait for Clk_period;
		Addr <=  "0001001011111";
		Trees_din <= x"0a01f708";
		wait for Clk_period;
		Addr <=  "0001001100000";
		Trees_din <= x"0d006704";
		wait for Clk_period;
		Addr <=  "0001001100001";
		Trees_din <= x"009e09e1";
		wait for Clk_period;
		Addr <=  "0001001100010";
		Trees_din <= x"ffa309e1";
		wait for Clk_period;
		Addr <=  "0001001100011";
		Trees_din <= x"ff5f09e1";
		wait for Clk_period;
		Addr <=  "0001001100100";
		Trees_din <= x"0605df08";
		wait for Clk_period;
		Addr <=  "0001001100101";
		Trees_din <= x"03fe2504";
		wait for Clk_period;
		Addr <=  "0001001100110";
		Trees_din <= x"00ba09e1";
		wait for Clk_period;
		Addr <=  "0001001100111";
		Trees_din <= x"005209e1";
		wait for Clk_period;
		Addr <=  "0001001101000";
		Trees_din <= x"0b00ac04";
		wait for Clk_period;
		Addr <=  "0001001101001";
		Trees_din <= x"ff6b09e1";
		wait for Clk_period;
		Addr <=  "0001001101010";
		Trees_din <= x"008909e1";
		wait for Clk_period;
		Addr <=  "0001001101011";
		Trees_din <= x"1b028110";
		wait for Clk_period;
		Addr <=  "0001001101100";
		Trees_din <= x"0e002108";
		wait for Clk_period;
		Addr <=  "0001001101101";
		Trees_din <= x"0d008b04";
		wait for Clk_period;
		Addr <=  "0001001101110";
		Trees_din <= x"ff4209e1";
		wait for Clk_period;
		Addr <=  "0001001101111";
		Trees_din <= x"009209e1";
		wait for Clk_period;
		Addr <=  "0001001110000";
		Trees_din <= x"02fda004";
		wait for Clk_period;
		Addr <=  "0001001110001";
		Trees_din <= x"00ac09e1";
		wait for Clk_period;
		Addr <=  "0001001110010";
		Trees_din <= x"ff8a09e1";
		wait for Clk_period;
		Addr <=  "0001001110011";
		Trees_din <= x"06f8e108";
		wait for Clk_period;
		Addr <=  "0001001110100";
		Trees_din <= x"1c028504";
		wait for Clk_period;
		Addr <=  "0001001110101";
		Trees_din <= x"fffc09e1";
		wait for Clk_period;
		Addr <=  "0001001110110";
		Trees_din <= x"007609e1";
		wait for Clk_period;
		Addr <=  "0001001110111";
		Trees_din <= x"ff0b09e1";
		wait for Clk_period;
		Addr <=  "0001001111000";
		Trees_din <= x"04042e60";
		wait for Clk_period;
		Addr <=  "0001001111001";
		Trees_din <= x"0400c424";
		wait for Clk_period;
		Addr <=  "0001001111010";
		Trees_din <= x"08004114";
		wait for Clk_period;
		Addr <=  "0001001111011";
		Trees_din <= x"1b026610";
		wait for Clk_period;
		Addr <=  "0001001111100";
		Trees_din <= x"1d025c08";
		wait for Clk_period;
		Addr <=  "0001001111101";
		Trees_din <= x"1501b204";
		wait for Clk_period;
		Addr <=  "0001001111110";
		Trees_din <= x"ff790b55";
		wait for Clk_period;
		Addr <=  "0001001111111";
		Trees_din <= x"002d0b55";
		wait for Clk_period;
		Addr <=  "0001010000000";
		Trees_din <= x"00fe5a04";
		wait for Clk_period;
		Addr <=  "0001010000001";
		Trees_din <= x"020f0b55";
		wait for Clk_period;
		Addr <=  "0001010000010";
		Trees_din <= x"00010b55";
		wait for Clk_period;
		Addr <=  "0001010000011";
		Trees_din <= x"ff6c0b55";
		wait for Clk_period;
		Addr <=  "0001010000100";
		Trees_din <= x"09002204";
		wait for Clk_period;
		Addr <=  "0001010000101";
		Trees_din <= x"00250b55";
		wait for Clk_period;
		Addr <=  "0001010000110";
		Trees_din <= x"09004d04";
		wait for Clk_period;
		Addr <=  "0001010000111";
		Trees_din <= x"ff650b55";
		wait for Clk_period;
		Addr <=  "0001010001000";
		Trees_din <= x"1603eb04";
		wait for Clk_period;
		Addr <=  "0001010001001";
		Trees_din <= x"ff9e0b55";
		wait for Clk_period;
		Addr <=  "0001010001010";
		Trees_din <= x"00400b55";
		wait for Clk_period;
		Addr <=  "0001010001011";
		Trees_din <= x"03ffdb20";
		wait for Clk_period;
		Addr <=  "0001010001100";
		Trees_din <= x"0c02e210";
		wait for Clk_period;
		Addr <=  "0001010001101";
		Trees_din <= x"03fcf208";
		wait for Clk_period;
		Addr <=  "0001010001110";
		Trees_din <= x"07ff8904";
		wait for Clk_period;
		Addr <=  "0001010001111";
		Trees_din <= x"00780b55";
		wait for Clk_period;
		Addr <=  "0001010010000";
		Trees_din <= x"ffc60b55";
		wait for Clk_period;
		Addr <=  "0001010010001";
		Trees_din <= x"0b012704";
		wait for Clk_period;
		Addr <=  "0001010010010";
		Trees_din <= x"ff9e0b55";
		wait for Clk_period;
		Addr <=  "0001010010011";
		Trees_din <= x"00db0b55";
		wait for Clk_period;
		Addr <=  "0001010010100";
		Trees_din <= x"03fd3908";
		wait for Clk_period;
		Addr <=  "0001010010101";
		Trees_din <= x"14003d04";
		wait for Clk_period;
		Addr <=  "0001010010110";
		Trees_din <= x"00270b55";
		wait for Clk_period;
		Addr <=  "0001010010111";
		Trees_din <= x"ff800b55";
		wait for Clk_period;
		Addr <=  "0001010011000";
		Trees_din <= x"0b00e704";
		wait for Clk_period;
		Addr <=  "0001010011001";
		Trees_din <= x"00e80b55";
		wait for Clk_period;
		Addr <=  "0001010011010";
		Trees_din <= x"ff950b55";
		wait for Clk_period;
		Addr <=  "0001010011011";
		Trees_din <= x"1300bc10";
		wait for Clk_period;
		Addr <=  "0001010011100";
		Trees_din <= x"15f78808";
		wait for Clk_period;
		Addr <=  "0001010011101";
		Trees_din <= x"0402e704";
		wait for Clk_period;
		Addr <=  "0001010011110";
		Trees_din <= x"fffd0b55";
		wait for Clk_period;
		Addr <=  "0001010011111";
		Trees_din <= x"00da0b55";
		wait for Clk_period;
		Addr <=  "0001010100000";
		Trees_din <= x"1afb5304";
		wait for Clk_period;
		Addr <=  "0001010100001";
		Trees_din <= x"00340b55";
		wait for Clk_period;
		Addr <=  "0001010100010";
		Trees_din <= x"ff8d0b55";
		wait for Clk_period;
		Addr <=  "0001010100011";
		Trees_din <= x"12003304";
		wait for Clk_period;
		Addr <=  "0001010100100";
		Trees_din <= x"ff790b55";
		wait for Clk_period;
		Addr <=  "0001010100101";
		Trees_din <= x"0403a504";
		wait for Clk_period;
		Addr <=  "0001010100110";
		Trees_din <= x"00f70b55";
		wait for Clk_period;
		Addr <=  "0001010100111";
		Trees_din <= x"ff980b55";
		wait for Clk_period;
		Addr <=  "0001010101000";
		Trees_din <= x"04095324";
		wait for Clk_period;
		Addr <=  "0001010101001";
		Trees_din <= x"00031a20";
		wait for Clk_period;
		Addr <=  "0001010101010";
		Trees_din <= x"01fff110";
		wait for Clk_period;
		Addr <=  "0001010101011";
		Trees_din <= x"12005c08";
		wait for Clk_period;
		Addr <=  "0001010101100";
		Trees_din <= x"13006904";
		wait for Clk_period;
		Addr <=  "0001010101101";
		Trees_din <= x"00a80b55";
		wait for Clk_period;
		Addr <=  "0001010101110";
		Trees_din <= x"003b0b55";
		wait for Clk_period;
		Addr <=  "0001010101111";
		Trees_din <= x"04069004";
		wait for Clk_period;
		Addr <=  "0001010110000";
		Trees_din <= x"ff5a0b55";
		wait for Clk_period;
		Addr <=  "0001010110001";
		Trees_din <= x"00330b55";
		wait for Clk_period;
		Addr <=  "0001010110010";
		Trees_din <= x"12003c08";
		wait for Clk_period;
		Addr <=  "0001010110011";
		Trees_din <= x"1afc3504";
		wait for Clk_period;
		Addr <=  "0001010110100";
		Trees_din <= x"ffbd0b55";
		wait for Clk_period;
		Addr <=  "0001010110101";
		Trees_din <= x"00e20b55";
		wait for Clk_period;
		Addr <=  "0001010110110";
		Trees_din <= x"05fbe904";
		wait for Clk_period;
		Addr <=  "0001010110111";
		Trees_din <= x"00630b55";
		wait for Clk_period;
		Addr <=  "0001010111000";
		Trees_din <= x"ff6a0b55";
		wait for Clk_period;
		Addr <=  "0001010111001";
		Trees_din <= x"ff750b55";
		wait for Clk_period;
		Addr <=  "0001010111010";
		Trees_din <= x"0705d220";
		wait for Clk_period;
		Addr <=  "0001010111011";
		Trees_din <= x"02fe2f10";
		wait for Clk_period;
		Addr <=  "0001010111100";
		Trees_din <= x"0a022108";
		wait for Clk_period;
		Addr <=  "0001010111101";
		Trees_din <= x"0101b404";
		wait for Clk_period;
		Addr <=  "0001010111110";
		Trees_din <= x"00a10b55";
		wait for Clk_period;
		Addr <=  "0001010111111";
		Trees_din <= x"00140b55";
		wait for Clk_period;
		Addr <=  "0001011000000";
		Trees_din <= x"1000f104";
		wait for Clk_period;
		Addr <=  "0001011000001";
		Trees_din <= x"ff1d0b55";
		wait for Clk_period;
		Addr <=  "0001011000010";
		Trees_din <= x"00710b55";
		wait for Clk_period;
		Addr <=  "0001011000011";
		Trees_din <= x"040d9708";
		wait for Clk_period;
		Addr <=  "0001011000100";
		Trees_din <= x"19000104";
		wait for Clk_period;
		Addr <=  "0001011000101";
		Trees_din <= x"ff650b55";
		wait for Clk_period;
		Addr <=  "0001011000110";
		Trees_din <= x"006c0b55";
		wait for Clk_period;
		Addr <=  "0001011000111";
		Trees_din <= x"09004404";
		wait for Clk_period;
		Addr <=  "0001011001000";
		Trees_din <= x"00a70b55";
		wait for Clk_period;
		Addr <=  "0001011001001";
		Trees_din <= x"00210b55";
		wait for Clk_period;
		Addr <=  "0001011001010";
		Trees_din <= x"040b000c";
		wait for Clk_period;
		Addr <=  "0001011001011";
		Trees_din <= x"0a00e304";
		wait for Clk_period;
		Addr <=  "0001011001100";
		Trees_din <= x"ff520b55";
		wait for Clk_period;
		Addr <=  "0001011001101";
		Trees_din <= x"05fd0104";
		wait for Clk_period;
		Addr <=  "0001011001110";
		Trees_din <= x"00800b55";
		wait for Clk_period;
		Addr <=  "0001011001111";
		Trees_din <= x"ff9d0b55";
		wait for Clk_period;
		Addr <=  "0001011010000";
		Trees_din <= x"16030304";
		wait for Clk_period;
		Addr <=  "0001011010001";
		Trees_din <= x"ffbd0b55";
		wait for Clk_period;
		Addr <=  "0001011010010";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "0001011010011";
		Trees_din <= x"ffc50b55";
		wait for Clk_period;
		Addr <=  "0001011010100";
		Trees_din <= x"00bc0b55";
		wait for Clk_period;
		Addr <=  "0001011010101";
		Trees_din <= x"0403332c";
		wait for Clk_period;
		Addr <=  "0001011010110";
		Trees_din <= x"04fb9604";
		wait for Clk_period;
		Addr <=  "0001011010111";
		Trees_din <= x"ff690c41";
		wait for Clk_period;
		Addr <=  "0001011011000";
		Trees_din <= x"1800841c";
		wait for Clk_period;
		Addr <=  "0001011011001";
		Trees_din <= x"060c0f10";
		wait for Clk_period;
		Addr <=  "0001011011010";
		Trees_din <= x"060b5f08";
		wait for Clk_period;
		Addr <=  "0001011011011";
		Trees_din <= x"1b026404";
		wait for Clk_period;
		Addr <=  "0001011011100";
		Trees_din <= x"003a0c41";
		wait for Clk_period;
		Addr <=  "0001011011101";
		Trees_din <= x"ffc20c41";
		wait for Clk_period;
		Addr <=  "0001011011110";
		Trees_din <= x"05fea704";
		wait for Clk_period;
		Addr <=  "0001011011111";
		Trees_din <= x"ffdf0c41";
		wait for Clk_period;
		Addr <=  "0001011100000";
		Trees_din <= x"01c10c41";
		wait for Clk_period;
		Addr <=  "0001011100001";
		Trees_din <= x"08003a04";
		wait for Clk_period;
		Addr <=  "0001011100010";
		Trees_din <= x"00aa0c41";
		wait for Clk_period;
		Addr <=  "0001011100011";
		Trees_din <= x"0b006804";
		wait for Clk_period;
		Addr <=  "0001011100100";
		Trees_din <= x"00530c41";
		wait for Clk_period;
		Addr <=  "0001011100101";
		Trees_din <= x"ff690c41";
		wait for Clk_period;
		Addr <=  "0001011100110";
		Trees_din <= x"18009a04";
		wait for Clk_period;
		Addr <=  "0001011100111";
		Trees_din <= x"ff640c41";
		wait for Clk_period;
		Addr <=  "0001011101000";
		Trees_din <= x"13006b04";
		wait for Clk_period;
		Addr <=  "0001011101001";
		Trees_din <= x"ff970c41";
		wait for Clk_period;
		Addr <=  "0001011101010";
		Trees_din <= x"009e0c41";
		wait for Clk_period;
		Addr <=  "0001011101011";
		Trees_din <= x"040b2b34";
		wait for Clk_period;
		Addr <=  "0001011101100";
		Trees_din <= x"04068420";
		wait for Clk_period;
		Addr <=  "0001011101101";
		Trees_din <= x"07ff9810";
		wait for Clk_period;
		Addr <=  "0001011101110";
		Trees_din <= x"11000008";
		wait for Clk_period;
		Addr <=  "0001011101111";
		Trees_din <= x"17040004";
		wait for Clk_period;
		Addr <=  "0001011110000";
		Trees_din <= x"011f0c41";
		wait for Clk_period;
		Addr <=  "0001011110001";
		Trees_din <= x"00080c41";
		wait for Clk_period;
		Addr <=  "0001011110010";
		Trees_din <= x"060c0004";
		wait for Clk_period;
		Addr <=  "0001011110011";
		Trees_din <= x"00380c41";
		wait for Clk_period;
		Addr <=  "0001011110100";
		Trees_din <= x"ff870c41";
		wait for Clk_period;
		Addr <=  "0001011110101";
		Trees_din <= x"05ff3c08";
		wait for Clk_period;
		Addr <=  "0001011110110";
		Trees_din <= x"0e003604";
		wait for Clk_period;
		Addr <=  "0001011110111";
		Trees_din <= x"ffe10c41";
		wait for Clk_period;
		Addr <=  "0001011111000";
		Trees_din <= x"00360c41";
		wait for Clk_period;
		Addr <=  "0001011111001";
		Trees_din <= x"05ff7504";
		wait for Clk_period;
		Addr <=  "0001011111010";
		Trees_din <= x"01570c41";
		wait for Clk_period;
		Addr <=  "0001011111011";
		Trees_din <= x"00350c41";
		wait for Clk_period;
		Addr <=  "0001011111100";
		Trees_din <= x"0101b410";
		wait for Clk_period;
		Addr <=  "0001011111101";
		Trees_din <= x"19000208";
		wait for Clk_period;
		Addr <=  "0001011111110";
		Trees_din <= x"1703d604";
		wait for Clk_period;
		Addr <=  "0001011111111";
		Trees_din <= x"00150c41";
		wait for Clk_period;
		Addr <=  "0001100000000";
		Trees_din <= x"00570c41";
		wait for Clk_period;
		Addr <=  "0001100000001";
		Trees_din <= x"1703e504";
		wait for Clk_period;
		Addr <=  "0001100000010";
		Trees_din <= x"007d0c41";
		wait for Clk_period;
		Addr <=  "0001100000011";
		Trees_din <= x"000b0c41";
		wait for Clk_period;
		Addr <=  "0001100000100";
		Trees_din <= x"ff650c41";
		wait for Clk_period;
		Addr <=  "0001100000101";
		Trees_din <= x"0003ad14";
		wait for Clk_period;
		Addr <=  "0001100000110";
		Trees_din <= x"1600d108";
		wait for Clk_period;
		Addr <=  "0001100000111";
		Trees_din <= x"02fb5f04";
		wait for Clk_period;
		Addr <=  "0001100001000";
		Trees_din <= x"ffa10c41";
		wait for Clk_period;
		Addr <=  "0001100001001";
		Trees_din <= x"006b0c41";
		wait for Clk_period;
		Addr <=  "0001100001010";
		Trees_din <= x"07fb7f04";
		wait for Clk_period;
		Addr <=  "0001100001011";
		Trees_din <= x"fffd0c41";
		wait for Clk_period;
		Addr <=  "0001100001100";
		Trees_din <= x"21000b04";
		wait for Clk_period;
		Addr <=  "0001100001101";
		Trees_din <= x"009e0c41";
		wait for Clk_period;
		Addr <=  "0001100001110";
		Trees_din <= x"001a0c41";
		wait for Clk_period;
		Addr <=  "0001100001111";
		Trees_din <= x"ffe10c41";
		wait for Clk_period;
		Addr <=  "0001100010000";
		Trees_din <= x"0401d230";
		wait for Clk_period;
		Addr <=  "0001100010001";
		Trees_din <= x"1b026618";
		wait for Clk_period;
		Addr <=  "0001100010010";
		Trees_din <= x"1afc6704";
		wait for Clk_period;
		Addr <=  "0001100010011";
		Trees_din <= x"01520d35";
		wait for Clk_period;
		Addr <=  "0001100010100";
		Trees_din <= x"09004a10";
		wait for Clk_period;
		Addr <=  "0001100010101";
		Trees_din <= x"0f007308";
		wait for Clk_period;
		Addr <=  "0001100010110";
		Trees_din <= x"0c018504";
		wait for Clk_period;
		Addr <=  "0001100010111";
		Trees_din <= x"ffce0d35";
		wait for Clk_period;
		Addr <=  "0001100011000";
		Trees_din <= x"00cd0d35";
		wait for Clk_period;
		Addr <=  "0001100011001";
		Trees_din <= x"1ffd6204";
		wait for Clk_period;
		Addr <=  "0001100011010";
		Trees_din <= x"ffef0d35";
		wait for Clk_period;
		Addr <=  "0001100011011";
		Trees_din <= x"ff6b0d35";
		wait for Clk_period;
		Addr <=  "0001100011100";
		Trees_din <= x"00c90d35";
		wait for Clk_period;
		Addr <=  "0001100011101";
		Trees_din <= x"19008310";
		wait for Clk_period;
		Addr <=  "0001100011110";
		Trees_din <= x"09004c08";
		wait for Clk_period;
		Addr <=  "0001100011111";
		Trees_din <= x"00fba204";
		wait for Clk_period;
		Addr <=  "0001100100000";
		Trees_din <= x"00360d35";
		wait for Clk_period;
		Addr <=  "0001100100001";
		Trees_din <= x"ff660d35";
		wait for Clk_period;
		Addr <=  "0001100100010";
		Trees_din <= x"0c027104";
		wait for Clk_period;
		Addr <=  "0001100100011";
		Trees_din <= x"ff8c0d35";
		wait for Clk_period;
		Addr <=  "0001100100100";
		Trees_din <= x"009b0d35";
		wait for Clk_period;
		Addr <=  "0001100100101";
		Trees_din <= x"07fe6404";
		wait for Clk_period;
		Addr <=  "0001100100110";
		Trees_din <= x"ffad0d35";
		wait for Clk_period;
		Addr <=  "0001100100111";
		Trees_din <= x"00d10d35";
		wait for Clk_period;
		Addr <=  "0001100101000";
		Trees_din <= x"040b2b28";
		wait for Clk_period;
		Addr <=  "0001100101001";
		Trees_din <= x"00031a20";
		wait for Clk_period;
		Addr <=  "0001100101010";
		Trees_din <= x"04056710";
		wait for Clk_period;
		Addr <=  "0001100101011";
		Trees_din <= x"02fb1f08";
		wait for Clk_period;
		Addr <=  "0001100101100";
		Trees_din <= x"09004c04";
		wait for Clk_period;
		Addr <=  "0001100101101";
		Trees_din <= x"ffe40d35";
		wait for Clk_period;
		Addr <=  "0001100101110";
		Trees_din <= x"00b60d35";
		wait for Clk_period;
		Addr <=  "0001100101111";
		Trees_din <= x"02fb2a04";
		wait for Clk_period;
		Addr <=  "0001100110000";
		Trees_din <= x"01300d35";
		wait for Clk_period;
		Addr <=  "0001100110001";
		Trees_din <= x"00210d35";
		wait for Clk_period;
		Addr <=  "0001100110010";
		Trees_din <= x"01fff108";
		wait for Clk_period;
		Addr <=  "0001100110011";
		Trees_din <= x"07001f04";
		wait for Clk_period;
		Addr <=  "0001100110100";
		Trees_din <= x"004b0d35";
		wait for Clk_period;
		Addr <=  "0001100110101";
		Trees_din <= x"00250d35";
		wait for Clk_period;
		Addr <=  "0001100110110";
		Trees_din <= x"05fca004";
		wait for Clk_period;
		Addr <=  "0001100110111";
		Trees_din <= x"00480d35";
		wait for Clk_period;
		Addr <=  "0001100111000";
		Trees_din <= x"ff980d35";
		wait for Clk_period;
		Addr <=  "0001100111001";
		Trees_din <= x"1300ca04";
		wait for Clk_period;
		Addr <=  "0001100111010";
		Trees_din <= x"ff700d35";
		wait for Clk_period;
		Addr <=  "0001100111011";
		Trees_din <= x"ffea0d35";
		wait for Clk_period;
		Addr <=  "0001100111100";
		Trees_din <= x"05fd2e0c";
		wait for Clk_period;
		Addr <=  "0001100111101";
		Trees_din <= x"0a022804";
		wait for Clk_period;
		Addr <=  "0001100111110";
		Trees_din <= x"00a80d35";
		wait for Clk_period;
		Addr <=  "0001100111111";
		Trees_din <= x"0b00b904";
		wait for Clk_period;
		Addr <=  "0001101000000";
		Trees_din <= x"00640d35";
		wait for Clk_period;
		Addr <=  "0001101000001";
		Trees_din <= x"ff910d35";
		wait for Clk_period;
		Addr <=  "0001101000010";
		Trees_din <= x"040e5410";
		wait for Clk_period;
		Addr <=  "0001101000011";
		Trees_din <= x"01006308";
		wait for Clk_period;
		Addr <=  "0001101000100";
		Trees_din <= x"18005604";
		wait for Clk_period;
		Addr <=  "0001101000101";
		Trees_din <= x"ffd90d35";
		wait for Clk_period;
		Addr <=  "0001101000110";
		Trees_din <= x"00910d35";
		wait for Clk_period;
		Addr <=  "0001101000111";
		Trees_din <= x"03fc4104";
		wait for Clk_period;
		Addr <=  "0001101001000";
		Trees_din <= x"ff360d35";
		wait for Clk_period;
		Addr <=  "0001101001001";
		Trees_din <= x"00220d35";
		wait for Clk_period;
		Addr <=  "0001101001010";
		Trees_din <= x"00facd04";
		wait for Clk_period;
		Addr <=  "0001101001011";
		Trees_din <= x"00070d35";
		wait for Clk_period;
		Addr <=  "0001101001100";
		Trees_din <= x"00a60d35";
		wait for Clk_period;
		Addr <=  "0001101001101";
		Trees_din <= x"0401c428";
		wait for Clk_period;
		Addr <=  "0001101001110";
		Trees_din <= x"04fb9604";
		wait for Clk_period;
		Addr <=  "0001101001111";
		Trees_din <= x"ff6d0df9";
		wait for Clk_period;
		Addr <=  "0001101010000";
		Trees_din <= x"03004a04";
		wait for Clk_period;
		Addr <=  "0001101010001";
		Trees_din <= x"ff6c0df9";
		wait for Clk_period;
		Addr <=  "0001101010010";
		Trees_din <= x"1b026610";
		wait for Clk_period;
		Addr <=  "0001101010011";
		Trees_din <= x"1d025e08";
		wait for Clk_period;
		Addr <=  "0001101010100";
		Trees_din <= x"0b00f704";
		wait for Clk_period;
		Addr <=  "0001101010101";
		Trees_din <= x"ffba0df9";
		wait for Clk_period;
		Addr <=  "0001101010110";
		Trees_din <= x"00d10df9";
		wait for Clk_period;
		Addr <=  "0001101010111";
		Trees_din <= x"08004104";
		wait for Clk_period;
		Addr <=  "0001101011000";
		Trees_din <= x"013f0df9";
		wait for Clk_period;
		Addr <=  "0001101011001";
		Trees_din <= x"00180df9";
		wait for Clk_period;
		Addr <=  "0001101011010";
		Trees_din <= x"1c028308";
		wait for Clk_period;
		Addr <=  "0001101011011";
		Trees_din <= x"0401a704";
		wait for Clk_period;
		Addr <=  "0001101011100";
		Trees_din <= x"ff700df9";
		wait for Clk_period;
		Addr <=  "0001101011101";
		Trees_din <= x"00320df9";
		wait for Clk_period;
		Addr <=  "0001101011110";
		Trees_din <= x"1300be04";
		wait for Clk_period;
		Addr <=  "0001101011111";
		Trees_din <= x"ff920df9";
		wait for Clk_period;
		Addr <=  "0001101100000";
		Trees_din <= x"00a30df9";
		wait for Clk_period;
		Addr <=  "0001101100001";
		Trees_din <= x"040b2b1c";
		wait for Clk_period;
		Addr <=  "0001101100010";
		Trees_din <= x"00031a14";
		wait for Clk_period;
		Addr <=  "0001101100011";
		Trees_din <= x"060d6810";
		wait for Clk_period;
		Addr <=  "0001101100100";
		Trees_din <= x"07019808";
		wait for Clk_period;
		Addr <=  "0001101100101";
		Trees_din <= x"09004204";
		wait for Clk_period;
		Addr <=  "0001101100110";
		Trees_din <= x"00390df9";
		wait for Clk_period;
		Addr <=  "0001101100111";
		Trees_din <= x"000e0df9";
		wait for Clk_period;
		Addr <=  "0001101101000";
		Trees_din <= x"06079a04";
		wait for Clk_period;
		Addr <=  "0001101101001";
		Trees_din <= x"00160df9";
		wait for Clk_period;
		Addr <=  "0001101101010";
		Trees_din <= x"ff8f0df9";
		wait for Clk_period;
		Addr <=  "0001101101011";
		Trees_din <= x"ff7c0df9";
		wait for Clk_period;
		Addr <=  "0001101101100";
		Trees_din <= x"1300cf04";
		wait for Clk_period;
		Addr <=  "0001101101101";
		Trees_din <= x"ff740df9";
		wait for Clk_period;
		Addr <=  "0001101101110";
		Trees_din <= x"ffec0df9";
		wait for Clk_period;
		Addr <=  "0001101101111";
		Trees_din <= x"05fd2e0c";
		wait for Clk_period;
		Addr <=  "0001101110000";
		Trees_din <= x"0a022804";
		wait for Clk_period;
		Addr <=  "0001101110001";
		Trees_din <= x"00a20df9";
		wait for Clk_period;
		Addr <=  "0001101110010";
		Trees_din <= x"0b00b904";
		wait for Clk_period;
		Addr <=  "0001101110011";
		Trees_din <= x"005d0df9";
		wait for Clk_period;
		Addr <=  "0001101110100";
		Trees_din <= x"ffa00df9";
		wait for Clk_period;
		Addr <=  "0001101110101";
		Trees_din <= x"05fd4204";
		wait for Clk_period;
		Addr <=  "0001101110110";
		Trees_din <= x"ff8b0df9";
		wait for Clk_period;
		Addr <=  "0001101110111";
		Trees_din <= x"0c000a08";
		wait for Clk_period;
		Addr <=  "0001101111000";
		Trees_din <= x"07032204";
		wait for Clk_period;
		Addr <=  "0001101111001";
		Trees_din <= x"00560df9";
		wait for Clk_period;
		Addr <=  "0001101111010";
		Trees_din <= x"ff6d0df9";
		wait for Clk_period;
		Addr <=  "0001101111011";
		Trees_din <= x"14004b04";
		wait for Clk_period;
		Addr <=  "0001101111100";
		Trees_din <= x"00910df9";
		wait for Clk_period;
		Addr <=  "0001101111101";
		Trees_din <= x"ffe20df9";
		wait for Clk_period;
		Addr <=  "0001101111110";
		Trees_din <= x"0400c424";
		wait for Clk_period;
		Addr <=  "0001101111111";
		Trees_din <= x"08004118";
		wait for Clk_period;
		Addr <=  "0001110000000";
		Trees_din <= x"1c026610";
		wait for Clk_period;
		Addr <=  "0001110000001";
		Trees_din <= x"1d025c04";
		wait for Clk_period;
		Addr <=  "0001110000010";
		Trees_din <= x"ff8f0efd";
		wait for Clk_period;
		Addr <=  "0001110000011";
		Trees_din <= x"0a00d008";
		wait for Clk_period;
		Addr <=  "0001110000100";
		Trees_din <= x"0a007404";
		wait for Clk_period;
		Addr <=  "0001110000101";
		Trees_din <= x"00410efd";
		wait for Clk_period;
		Addr <=  "0001110000110";
		Trees_din <= x"01bb0efd";
		wait for Clk_period;
		Addr <=  "0001110000111";
		Trees_din <= x"000c0efd";
		wait for Clk_period;
		Addr <=  "0001110001000";
		Trees_din <= x"1501b204";
		wait for Clk_period;
		Addr <=  "0001110001001";
		Trees_din <= x"ff770efd";
		wait for Clk_period;
		Addr <=  "0001110001010";
		Trees_din <= x"00290efd";
		wait for Clk_period;
		Addr <=  "0001110001011";
		Trees_din <= x"13005e04";
		wait for Clk_period;
		Addr <=  "0001110001100";
		Trees_din <= x"00420efd";
		wait for Clk_period;
		Addr <=  "0001110001101";
		Trees_din <= x"0b005404";
		wait for Clk_period;
		Addr <=  "0001110001110";
		Trees_din <= x"00080efd";
		wait for Clk_period;
		Addr <=  "0001110001111";
		Trees_din <= x"ff6a0efd";
		wait for Clk_period;
		Addr <=  "0001110010000";
		Trees_din <= x"04095330";
		wait for Clk_period;
		Addr <=  "0001110010001";
		Trees_din <= x"03fa4b10";
		wait for Clk_period;
		Addr <=  "0001110010010";
		Trees_din <= x"1300e10c";
		wait for Clk_period;
		Addr <=  "0001110010011";
		Trees_din <= x"00fd6704";
		wait for Clk_period;
		Addr <=  "0001110010100";
		Trees_din <= x"ff1b0efd";
		wait for Clk_period;
		Addr <=  "0001110010101";
		Trees_din <= x"04074204";
		wait for Clk_period;
		Addr <=  "0001110010110";
		Trees_din <= x"ff860efd";
		wait for Clk_period;
		Addr <=  "0001110010111";
		Trees_din <= x"002e0efd";
		wait for Clk_period;
		Addr <=  "0001110011000";
		Trees_din <= x"01000efd";
		wait for Clk_period;
		Addr <=  "0001110011001";
		Trees_din <= x"03fabd10";
		wait for Clk_period;
		Addr <=  "0001110011010";
		Trees_din <= x"08004108";
		wait for Clk_period;
		Addr <=  "0001110011011";
		Trees_din <= x"0e002a04";
		wait for Clk_period;
		Addr <=  "0001110011100";
		Trees_din <= x"ff650efd";
		wait for Clk_period;
		Addr <=  "0001110011101";
		Trees_din <= x"00360efd";
		wait for Clk_period;
		Addr <=  "0001110011110";
		Trees_din <= x"1e026704";
		wait for Clk_period;
		Addr <=  "0001110011111";
		Trees_din <= x"01010efd";
		wait for Clk_period;
		Addr <=  "0001110100000";
		Trees_din <= x"005c0efd";
		wait for Clk_period;
		Addr <=  "0001110100001";
		Trees_din <= x"05ff4708";
		wait for Clk_period;
		Addr <=  "0001110100010";
		Trees_din <= x"07ff7e04";
		wait for Clk_period;
		Addr <=  "0001110100011";
		Trees_din <= x"00260efd";
		wait for Clk_period;
		Addr <=  "0001110100100";
		Trees_din <= x"00030efd";
		wait for Clk_period;
		Addr <=  "0001110100101";
		Trees_din <= x"07fd9c04";
		wait for Clk_period;
		Addr <=  "0001110100110";
		Trees_din <= x"ffb90efd";
		wait for Clk_period;
		Addr <=  "0001110100111";
		Trees_din <= x"00680efd";
		wait for Clk_period;
		Addr <=  "0001110101000";
		Trees_din <= x"05fc2c18";
		wait for Clk_period;
		Addr <=  "0001110101001";
		Trees_din <= x"0704ef0c";
		wait for Clk_period;
		Addr <=  "0001110101010";
		Trees_din <= x"04096d04";
		wait for Clk_period;
		Addr <=  "0001110101011";
		Trees_din <= x"ffe60efd";
		wait for Clk_period;
		Addr <=  "0001110101100";
		Trees_din <= x"0f006504";
		wait for Clk_period;
		Addr <=  "0001110101101";
		Trees_din <= x"00190efd";
		wait for Clk_period;
		Addr <=  "0001110101110";
		Trees_din <= x"00a90efd";
		wait for Clk_period;
		Addr <=  "0001110101111";
		Trees_din <= x"0e002104";
		wait for Clk_period;
		Addr <=  "0001110110000";
		Trees_din <= x"ff7b0efd";
		wait for Clk_period;
		Addr <=  "0001110110001";
		Trees_din <= x"0b00b304";
		wait for Clk_period;
		Addr <=  "0001110110010";
		Trees_din <= x"ffe10efd";
		wait for Clk_period;
		Addr <=  "0001110110011";
		Trees_din <= x"00880efd";
		wait for Clk_period;
		Addr <=  "0001110110100";
		Trees_din <= x"040e5410";
		wait for Clk_period;
		Addr <=  "0001110110101";
		Trees_din <= x"01ffbf08";
		wait for Clk_period;
		Addr <=  "0001110110110";
		Trees_din <= x"0a022104";
		wait for Clk_period;
		Addr <=  "0001110110111";
		Trees_din <= x"00640efd";
		wait for Clk_period;
		Addr <=  "0001110111000";
		Trees_din <= x"ff880efd";
		wait for Clk_period;
		Addr <=  "0001110111001";
		Trees_din <= x"09003d04";
		wait for Clk_period;
		Addr <=  "0001110111010";
		Trees_din <= x"002a0efd";
		wait for Clk_period;
		Addr <=  "0001110111011";
		Trees_din <= x"ff860efd";
		wait for Clk_period;
		Addr <=  "0001110111100";
		Trees_din <= x"06d10d04";
		wait for Clk_period;
		Addr <=  "0001110111101";
		Trees_din <= x"00160efd";
		wait for Clk_period;
		Addr <=  "0001110111110";
		Trees_din <= x"009f0efd";
		wait for Clk_period;
		Addr <=  "0001110111111";
		Trees_din <= x"0400c424";
		wait for Clk_period;
		Addr <=  "0001111000000";
		Trees_din <= x"08004118";
		wait for Clk_period;
		Addr <=  "0001111000001";
		Trees_din <= x"1c026610";
		wait for Clk_period;
		Addr <=  "0001111000010";
		Trees_din <= x"1d025c04";
		wait for Clk_period;
		Addr <=  "0001111000011";
		Trees_din <= x"ff941001";
		wait for Clk_period;
		Addr <=  "0001111000100";
		Trees_din <= x"00fe5a08";
		wait for Clk_period;
		Addr <=  "0001111000101";
		Trees_din <= x"19000004";
		wait for Clk_period;
		Addr <=  "0001111000110";
		Trees_din <= x"00461001";
		wait for Clk_period;
		Addr <=  "0001111000111";
		Trees_din <= x"014a1001";
		wait for Clk_period;
		Addr <=  "0001111001000";
		Trees_din <= x"00111001";
		wait for Clk_period;
		Addr <=  "0001111001001";
		Trees_din <= x"13009704";
		wait for Clk_period;
		Addr <=  "0001111001010";
		Trees_din <= x"00221001";
		wait for Clk_period;
		Addr <=  "0001111001011";
		Trees_din <= x"ff7a1001";
		wait for Clk_period;
		Addr <=  "0001111001100";
		Trees_din <= x"13005e04";
		wait for Clk_period;
		Addr <=  "0001111001101";
		Trees_din <= x"003f1001";
		wait for Clk_period;
		Addr <=  "0001111001110";
		Trees_din <= x"00066304";
		wait for Clk_period;
		Addr <=  "0001111001111";
		Trees_din <= x"ff6b1001";
		wait for Clk_period;
		Addr <=  "0001111010000";
		Trees_din <= x"000f1001";
		wait for Clk_period;
		Addr <=  "0001111010001";
		Trees_din <= x"040b2b3c";
		wait for Clk_period;
		Addr <=  "0001111010010";
		Trees_din <= x"0b004b1c";
		wait for Clk_period;
		Addr <=  "0001111010011";
		Trees_din <= x"0900440c";
		wait for Clk_period;
		Addr <=  "0001111010100";
		Trees_din <= x"00fd4004";
		wait for Clk_period;
		Addr <=  "0001111010101";
		Trees_din <= x"ffe51001";
		wait for Clk_period;
		Addr <=  "0001111010110";
		Trees_din <= x"0d00ae04";
		wait for Clk_period;
		Addr <=  "0001111010111";
		Trees_din <= x"013f1001";
		wait for Clk_period;
		Addr <=  "0001111011000";
		Trees_din <= x"00661001";
		wait for Clk_period;
		Addr <=  "0001111011001";
		Trees_din <= x"04055c08";
		wait for Clk_period;
		Addr <=  "0001111011010";
		Trees_din <= x"15f81704";
		wait for Clk_period;
		Addr <=  "0001111011011";
		Trees_din <= x"00791001";
		wait for Clk_period;
		Addr <=  "0001111011100";
		Trees_din <= x"ff721001";
		wait for Clk_period;
		Addr <=  "0001111011101";
		Trees_din <= x"19000004";
		wait for Clk_period;
		Addr <=  "0001111011110";
		Trees_din <= x"ffba1001";
		wait for Clk_period;
		Addr <=  "0001111011111";
		Trees_din <= x"00b21001";
		wait for Clk_period;
		Addr <=  "0001111100000";
		Trees_din <= x"01ff8010";
		wait for Clk_period;
		Addr <=  "0001111100001";
		Trees_din <= x"1cfbec08";
		wait for Clk_period;
		Addr <=  "0001111100010";
		Trees_din <= x"0609e504";
		wait for Clk_period;
		Addr <=  "0001111100011";
		Trees_din <= x"ff7f1001";
		wait for Clk_period;
		Addr <=  "0001111100100";
		Trees_din <= x"003e1001";
		wait for Clk_period;
		Addr <=  "0001111100101";
		Trees_din <= x"0b00f904";
		wait for Clk_period;
		Addr <=  "0001111100110";
		Trees_din <= x"00141001";
		wait for Clk_period;
		Addr <=  "0001111100111";
		Trees_din <= x"00551001";
		wait for Clk_period;
		Addr <=  "0001111101000";
		Trees_din <= x"15f87008";
		wait for Clk_period;
		Addr <=  "0001111101001";
		Trees_din <= x"11001704";
		wait for Clk_period;
		Addr <=  "0001111101010";
		Trees_din <= x"ffd91001";
		wait for Clk_period;
		Addr <=  "0001111101011";
		Trees_din <= x"ff461001";
		wait for Clk_period;
		Addr <=  "0001111101100";
		Trees_din <= x"0f007404";
		wait for Clk_period;
		Addr <=  "0001111101101";
		Trees_din <= x"009c1001";
		wait for Clk_period;
		Addr <=  "0001111101110";
		Trees_din <= x"ffe91001";
		wait for Clk_period;
		Addr <=  "0001111101111";
		Trees_din <= x"05fd2e0c";
		wait for Clk_period;
		Addr <=  "0001111110000";
		Trees_din <= x"0e004908";
		wait for Clk_period;
		Addr <=  "0001111110001";
		Trees_din <= x"07079b04";
		wait for Clk_period;
		Addr <=  "0001111110010";
		Trees_din <= x"009c1001";
		wait for Clk_period;
		Addr <=  "0001111110011";
		Trees_din <= x"001f1001";
		wait for Clk_period;
		Addr <=  "0001111110100";
		Trees_din <= x"fffe1001";
		wait for Clk_period;
		Addr <=  "0001111110101";
		Trees_din <= x"040e5410";
		wait for Clk_period;
		Addr <=  "0001111110110";
		Trees_din <= x"01006308";
		wait for Clk_period;
		Addr <=  "0001111110111";
		Trees_din <= x"12003e04";
		wait for Clk_period;
		Addr <=  "0001111111000";
		Trees_din <= x"ffe71001";
		wait for Clk_period;
		Addr <=  "0001111111001";
		Trees_din <= x"007b1001";
		wait for Clk_period;
		Addr <=  "0001111111010";
		Trees_din <= x"03fc4104";
		wait for Clk_period;
		Addr <=  "0001111111011";
		Trees_din <= x"ff531001";
		wait for Clk_period;
		Addr <=  "0001111111100";
		Trees_din <= x"001b1001";
		wait for Clk_period;
		Addr <=  "0001111111101";
		Trees_din <= x"00facd04";
		wait for Clk_period;
		Addr <=  "0001111111110";
		Trees_din <= x"fffe1001";
		wait for Clk_period;
		Addr <=  "0001111111111";
		Trees_din <= x"00941001";
		wait for Clk_period;
		Addr <=  "0010000000000";
		Trees_din <= x"04fb9604";
		wait for Clk_period;
		Addr <=  "0010000000001";
		Trees_din <= x"ff741095";
		wait for Clk_period;
		Addr <=  "0010000000010";
		Trees_din <= x"040b2b24";
		wait for Clk_period;
		Addr <=  "0010000000011";
		Trees_din <= x"060d6820";
		wait for Clk_period;
		Addr <=  "0010000000100";
		Trees_din <= x"0700ca10";
		wait for Clk_period;
		Addr <=  "0010000000101";
		Trees_din <= x"18007f08";
		wait for Clk_period;
		Addr <=  "0010000000110";
		Trees_din <= x"18007c04";
		wait for Clk_period;
		Addr <=  "0010000000111";
		Trees_din <= x"001f1095";
		wait for Clk_period;
		Addr <=  "0010000001000";
		Trees_din <= x"00b81095";
		wait for Clk_period;
		Addr <=  "0010000001001";
		Trees_din <= x"05fd2e04";
		wait for Clk_period;
		Addr <=  "0010000001010";
		Trees_din <= x"00411095";
		wait for Clk_period;
		Addr <=  "0010000001011";
		Trees_din <= x"ffd31095";
		wait for Clk_period;
		Addr <=  "0010000001100";
		Trees_din <= x"04026608";
		wait for Clk_period;
		Addr <=  "0010000001101";
		Trees_din <= x"15f70f04";
		wait for Clk_period;
		Addr <=  "0010000001110";
		Trees_din <= x"00371095";
		wait for Clk_period;
		Addr <=  "0010000001111";
		Trees_din <= x"ff6a1095";
		wait for Clk_period;
		Addr <=  "0010000010000";
		Trees_din <= x"19000404";
		wait for Clk_period;
		Addr <=  "0010000010001";
		Trees_din <= x"fff91095";
		wait for Clk_period;
		Addr <=  "0010000010010";
		Trees_din <= x"002e1095";
		wait for Clk_period;
		Addr <=  "0010000010011";
		Trees_din <= x"ff791095";
		wait for Clk_period;
		Addr <=  "0010000010100";
		Trees_din <= x"05fd2e0c";
		wait for Clk_period;
		Addr <=  "0010000010101";
		Trees_din <= x"0a022804";
		wait for Clk_period;
		Addr <=  "0010000010110";
		Trees_din <= x"00961095";
		wait for Clk_period;
		Addr <=  "0010000010111";
		Trees_din <= x"19000004";
		wait for Clk_period;
		Addr <=  "0010000011000";
		Trees_din <= x"ffc31095";
		wait for Clk_period;
		Addr <=  "0010000011001";
		Trees_din <= x"005d1095";
		wait for Clk_period;
		Addr <=  "0010000011010";
		Trees_din <= x"040e5410";
		wait for Clk_period;
		Addr <=  "0010000011011";
		Trees_din <= x"01006308";
		wait for Clk_period;
		Addr <=  "0010000011100";
		Trees_din <= x"12003e04";
		wait for Clk_period;
		Addr <=  "0010000011101";
		Trees_din <= x"ffe71095";
		wait for Clk_period;
		Addr <=  "0010000011110";
		Trees_din <= x"00741095";
		wait for Clk_period;
		Addr <=  "0010000011111";
		Trees_din <= x"03fc4104";
		wait for Clk_period;
		Addr <=  "0010000100000";
		Trees_din <= x"ff641095";
		wait for Clk_period;
		Addr <=  "0010000100001";
		Trees_din <= x"00151095";
		wait for Clk_period;
		Addr <=  "0010000100010";
		Trees_din <= x"00facd04";
		wait for Clk_period;
		Addr <=  "0010000100011";
		Trees_din <= x"00011095";
		wait for Clk_period;
		Addr <=  "0010000100100";
		Trees_din <= x"008e1095";
		wait for Clk_period;
		Addr <=  "0010000100101";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0010000100110";
		Trees_din <= x"04fb9604";
		wait for Clk_period;
		Addr <=  "0010000100111";
		Trees_din <= x"ff77111d";
		wait for Clk_period;
		Addr <=  "0010000101000";
		Trees_din <= x"040b2b24";
		wait for Clk_period;
		Addr <=  "0010000101001";
		Trees_din <= x"060d6820";
		wait for Clk_period;
		Addr <=  "0010000101010";
		Trees_din <= x"0d009310";
		wait for Clk_period;
		Addr <=  "0010000101011";
		Trees_din <= x"2003fe08";
		wait for Clk_period;
		Addr <=  "0010000101100";
		Trees_din <= x"02fc5b04";
		wait for Clk_period;
		Addr <=  "0010000101101";
		Trees_din <= x"ff5a111d";
		wait for Clk_period;
		Addr <=  "0010000101110";
		Trees_din <= x"0033111d";
		wait for Clk_period;
		Addr <=  "0010000101111";
		Trees_din <= x"00001f04";
		wait for Clk_period;
		Addr <=  "0010000110000";
		Trees_din <= x"0012111d";
		wait for Clk_period;
		Addr <=  "0010000110001";
		Trees_din <= x"ffde111d";
		wait for Clk_period;
		Addr <=  "0010000110010";
		Trees_din <= x"1c026108";
		wait for Clk_period;
		Addr <=  "0010000110011";
		Trees_din <= x"0c00ec04";
		wait for Clk_period;
		Addr <=  "0010000110100";
		Trees_din <= x"ff88111d";
		wait for Clk_period;
		Addr <=  "0010000110101";
		Trees_din <= x"0059111d";
		wait for Clk_period;
		Addr <=  "0010000110110";
		Trees_din <= x"12002e04";
		wait for Clk_period;
		Addr <=  "0010000110111";
		Trees_din <= x"ffc6111d";
		wait for Clk_period;
		Addr <=  "0010000111000";
		Trees_din <= x"0068111d";
		wait for Clk_period;
		Addr <=  "0010000111001";
		Trees_din <= x"ff7e111d";
		wait for Clk_period;
		Addr <=  "0010000111010";
		Trees_din <= x"05fd2e0c";
		wait for Clk_period;
		Addr <=  "0010000111011";
		Trees_din <= x"0e004908";
		wait for Clk_period;
		Addr <=  "0010000111100";
		Trees_din <= x"07079b04";
		wait for Clk_period;
		Addr <=  "0010000111101";
		Trees_din <= x"0096111d";
		wait for Clk_period;
		Addr <=  "0010000111110";
		Trees_din <= x"0019111d";
		wait for Clk_period;
		Addr <=  "0010000111111";
		Trees_din <= x"fffb111d";
		wait for Clk_period;
		Addr <=  "0010001000000";
		Trees_din <= x"05fd4204";
		wait for Clk_period;
		Addr <=  "0010001000001";
		Trees_din <= x"ff97111d";
		wait for Clk_period;
		Addr <=  "0010001000010";
		Trees_din <= x"0c000a04";
		wait for Clk_period;
		Addr <=  "0010001000011";
		Trees_din <= x"ffcc111d";
		wait for Clk_period;
		Addr <=  "0010001000100";
		Trees_din <= x"09004704";
		wait for Clk_period;
		Addr <=  "0010001000101";
		Trees_din <= x"0081111d";
		wait for Clk_period;
		Addr <=  "0010001000110";
		Trees_din <= x"fff3111d";
		wait for Clk_period;
		Addr <=  "0010001000111";
		Trees_din <= x"04fb9604";
		wait for Clk_period;
		Addr <=  "0010001001000";
		Trees_din <= x"ff7a11c1";
		wait for Clk_period;
		Addr <=  "0010001001001";
		Trees_din <= x"040b2b30";
		wait for Clk_period;
		Addr <=  "0010001001010";
		Trees_din <= x"1200611c";
		wait for Clk_period;
		Addr <=  "0010001001011";
		Trees_din <= x"0706c610";
		wait for Clk_period;
		Addr <=  "0010001001100";
		Trees_din <= x"1b028808";
		wait for Clk_period;
		Addr <=  "0010001001101";
		Trees_din <= x"0d009e04";
		wait for Clk_period;
		Addr <=  "0010001001110";
		Trees_din <= x"000e11c1";
		wait for Clk_period;
		Addr <=  "0010001001111";
		Trees_din <= x"005011c1";
		wait for Clk_period;
		Addr <=  "0010001010000";
		Trees_din <= x"00fe5004";
		wait for Clk_period;
		Addr <=  "0010001010001";
		Trees_din <= x"ff8411c1";
		wait for Clk_period;
		Addr <=  "0010001010010";
		Trees_din <= x"001d11c1";
		wait for Clk_period;
		Addr <=  "0010001010011";
		Trees_din <= x"16040008";
		wait for Clk_period;
		Addr <=  "0010001010100";
		Trees_din <= x"03fd5504";
		wait for Clk_period;
		Addr <=  "0010001010101";
		Trees_din <= x"ff6a11c1";
		wait for Clk_period;
		Addr <=  "0010001010110";
		Trees_din <= x"fffd11c1";
		wait for Clk_period;
		Addr <=  "0010001010111";
		Trees_din <= x"004c11c1";
		wait for Clk_period;
		Addr <=  "0010001011000";
		Trees_din <= x"00fe880c";
		wait for Clk_period;
		Addr <=  "0010001011001";
		Trees_din <= x"0b00c808";
		wait for Clk_period;
		Addr <=  "0010001011010";
		Trees_din <= x"05fdd804";
		wait for Clk_period;
		Addr <=  "0010001011011";
		Trees_din <= x"ff3c11c1";
		wait for Clk_period;
		Addr <=  "0010001011100";
		Trees_din <= x"ffca11c1";
		wait for Clk_period;
		Addr <=  "0010001011101";
		Trees_din <= x"fff711c1";
		wait for Clk_period;
		Addr <=  "0010001011110";
		Trees_din <= x"0d006b04";
		wait for Clk_period;
		Addr <=  "0010001011111";
		Trees_din <= x"007211c1";
		wait for Clk_period;
		Addr <=  "0010001100000";
		Trees_din <= x"ff9f11c1";
		wait for Clk_period;
		Addr <=  "0010001100001";
		Trees_din <= x"02fd8114";
		wait for Clk_period;
		Addr <=  "0010001100010";
		Trees_din <= x"1600d104";
		wait for Clk_period;
		Addr <=  "0010001100011";
		Trees_din <= x"ffd811c1";
		wait for Clk_period;
		Addr <=  "0010001100100";
		Trees_din <= x"15f71d08";
		wait for Clk_period;
		Addr <=  "0010001100101";
		Trees_din <= x"0e002704";
		wait for Clk_period;
		Addr <=  "0010001100110";
		Trees_din <= x"ffc111c1";
		wait for Clk_period;
		Addr <=  "0010001100111";
		Trees_din <= x"005f11c1";
		wait for Clk_period;
		Addr <=  "0010001101000";
		Trees_din <= x"17026a04";
		wait for Clk_period;
		Addr <=  "0010001101001";
		Trees_din <= x"002911c1";
		wait for Clk_period;
		Addr <=  "0010001101010";
		Trees_din <= x"009111c1";
		wait for Clk_period;
		Addr <=  "0010001101011";
		Trees_din <= x"00024008";
		wait for Clk_period;
		Addr <=  "0010001101100";
		Trees_din <= x"09004404";
		wait for Clk_period;
		Addr <=  "0010001101101";
		Trees_din <= x"007611c1";
		wait for Clk_period;
		Addr <=  "0010001101110";
		Trees_din <= x"ffed11c1";
		wait for Clk_period;
		Addr <=  "0010001101111";
		Trees_din <= x"ff9911c1";
		wait for Clk_period;
		Addr <=  "0010001110000";
		Trees_din <= x"02fd8174";
		wait for Clk_period;
		Addr <=  "0010001110001";
		Trees_din <= x"04095340";
		wait for Clk_period;
		Addr <=  "0010001110010";
		Trees_din <= x"07fedb20";
		wait for Clk_period;
		Addr <=  "0010001110011";
		Trees_din <= x"03fcb210";
		wait for Clk_period;
		Addr <=  "0010001110100";
		Trees_din <= x"00fe1108";
		wait for Clk_period;
		Addr <=  "0010001110101";
		Trees_din <= x"1b028104";
		wait for Clk_period;
		Addr <=  "0010001110110";
		Trees_din <= x"00a3130d";
		wait for Clk_period;
		Addr <=  "0010001110111";
		Trees_din <= x"ff9d130d";
		wait for Clk_period;
		Addr <=  "0010001111000";
		Trees_din <= x"02fc4704";
		wait for Clk_period;
		Addr <=  "0010001111001";
		Trees_din <= x"ffdf130d";
		wait for Clk_period;
		Addr <=  "0010001111010";
		Trees_din <= x"012a130d";
		wait for Clk_period;
		Addr <=  "0010001111011";
		Trees_din <= x"00ff3308";
		wait for Clk_period;
		Addr <=  "0010001111100";
		Trees_din <= x"0a007904";
		wait for Clk_period;
		Addr <=  "0010001111101";
		Trees_din <= x"ffca130d";
		wait for Clk_period;
		Addr <=  "0010001111110";
		Trees_din <= x"002b130d";
		wait for Clk_period;
		Addr <=  "0010001111111";
		Trees_din <= x"0a01c304";
		wait for Clk_period;
		Addr <=  "0010010000000";
		Trees_din <= x"0096130d";
		wait for Clk_period;
		Addr <=  "0010010000001";
		Trees_din <= x"ff6c130d";
		wait for Clk_period;
		Addr <=  "0010010000010";
		Trees_din <= x"0c02c510";
		wait for Clk_period;
		Addr <=  "0010010000011";
		Trees_din <= x"0a011b08";
		wait for Clk_period;
		Addr <=  "0010010000100";
		Trees_din <= x"1bfaf204";
		wait for Clk_period;
		Addr <=  "0010010000101";
		Trees_din <= x"ff97130d";
		wait for Clk_period;
		Addr <=  "0010010000110";
		Trees_din <= x"000d130d";
		wait for Clk_period;
		Addr <=  "0010010000111";
		Trees_din <= x"1e027904";
		wait for Clk_period;
		Addr <=  "0010010001000";
		Trees_din <= x"ffac130d";
		wait for Clk_period;
		Addr <=  "0010010001001";
		Trees_din <= x"0015130d";
		wait for Clk_period;
		Addr <=  "0010010001010";
		Trees_din <= x"1603f608";
		wait for Clk_period;
		Addr <=  "0010010001011";
		Trees_din <= x"0d006804";
		wait for Clk_period;
		Addr <=  "0010010001100";
		Trees_din <= x"ffc1130d";
		wait for Clk_period;
		Addr <=  "0010010001101";
		Trees_din <= x"008d130d";
		wait for Clk_period;
		Addr <=  "0010010001110";
		Trees_din <= x"0c02e204";
		wait for Clk_period;
		Addr <=  "0010010001111";
		Trees_din <= x"00b6130d";
		wait for Clk_period;
		Addr <=  "0010010010000";
		Trees_din <= x"ff47130d";
		wait for Clk_period;
		Addr <=  "0010010010001";
		Trees_din <= x"02fa5518";
		wait for Clk_period;
		Addr <=  "0010010010010";
		Trees_din <= x"0f00770c";
		wait for Clk_period;
		Addr <=  "0010010010011";
		Trees_din <= x"13008c08";
		wait for Clk_period;
		Addr <=  "0010010010100";
		Trees_din <= x"0f006b04";
		wait for Clk_period;
		Addr <=  "0010010010101";
		Trees_din <= x"0052130d";
		wait for Clk_period;
		Addr <=  "0010010010110";
		Trees_din <= x"ff88130d";
		wait for Clk_period;
		Addr <=  "0010010010111";
		Trees_din <= x"0092130d";
		wait for Clk_period;
		Addr <=  "0010010011000";
		Trees_din <= x"0f008808";
		wait for Clk_period;
		Addr <=  "0010010011001";
		Trees_din <= x"0c014004";
		wait for Clk_period;
		Addr <=  "0010010011010";
		Trees_din <= x"ff2e130d";
		wait for Clk_period;
		Addr <=  "0010010011011";
		Trees_din <= x"000d130d";
		wait for Clk_period;
		Addr <=  "0010010011100";
		Trees_din <= x"0068130d";
		wait for Clk_period;
		Addr <=  "0010010011101";
		Trees_din <= x"12004c0c";
		wait for Clk_period;
		Addr <=  "0010010011110";
		Trees_din <= x"0607db08";
		wait for Clk_period;
		Addr <=  "0010010011111";
		Trees_din <= x"1c023e04";
		wait for Clk_period;
		Addr <=  "0010010100000";
		Trees_din <= x"0011130d";
		wait for Clk_period;
		Addr <=  "0010010100001";
		Trees_din <= x"0095130d";
		wait for Clk_period;
		Addr <=  "0010010100010";
		Trees_din <= x"ffe9130d";
		wait for Clk_period;
		Addr <=  "0010010100011";
		Trees_din <= x"06026c08";
		wait for Clk_period;
		Addr <=  "0010010100100";
		Trees_din <= x"0601e804";
		wait for Clk_period;
		Addr <=  "0010010100101";
		Trees_din <= x"001c130d";
		wait for Clk_period;
		Addr <=  "0010010100110";
		Trees_din <= x"ff0a130d";
		wait for Clk_period;
		Addr <=  "0010010100111";
		Trees_din <= x"06038604";
		wait for Clk_period;
		Addr <=  "0010010101000";
		Trees_din <= x"0025130d";
		wait for Clk_period;
		Addr <=  "0010010101001";
		Trees_din <= x"0083130d";
		wait for Clk_period;
		Addr <=  "0010010101010";
		Trees_din <= x"0e00412c";
		wait for Clk_period;
		Addr <=  "0010010101011";
		Trees_din <= x"0d006610";
		wait for Clk_period;
		Addr <=  "0010010101100";
		Trees_din <= x"01fd9308";
		wait for Clk_period;
		Addr <=  "0010010101101";
		Trees_din <= x"13009604";
		wait for Clk_period;
		Addr <=  "0010010101110";
		Trees_din <= x"011d130d";
		wait for Clk_period;
		Addr <=  "0010010101111";
		Trees_din <= x"004e130d";
		wait for Clk_period;
		Addr <=  "0010010110000";
		Trees_din <= x"0a002f04";
		wait for Clk_period;
		Addr <=  "0010010110001";
		Trees_din <= x"0095130d";
		wait for Clk_period;
		Addr <=  "0010010110010";
		Trees_din <= x"ffae130d";
		wait for Clk_period;
		Addr <=  "0010010110011";
		Trees_din <= x"10022110";
		wait for Clk_period;
		Addr <=  "0010010110100";
		Trees_din <= x"1afd5908";
		wait for Clk_period;
		Addr <=  "0010010110101";
		Trees_din <= x"0c013104";
		wait for Clk_period;
		Addr <=  "0010010110110";
		Trees_din <= x"0013130d";
		wait for Clk_period;
		Addr <=  "0010010110111";
		Trees_din <= x"ffb1130d";
		wait for Clk_period;
		Addr <=  "0010010111000";
		Trees_din <= x"0e003104";
		wait for Clk_period;
		Addr <=  "0010010111001";
		Trees_din <= x"ff3b130d";
		wait for Clk_period;
		Addr <=  "0010010111010";
		Trees_din <= x"ffdb130d";
		wait for Clk_period;
		Addr <=  "0010010111011";
		Trees_din <= x"0d007604";
		wait for Clk_period;
		Addr <=  "0010010111100";
		Trees_din <= x"ff8a130d";
		wait for Clk_period;
		Addr <=  "0010010111101";
		Trees_din <= x"0e002404";
		wait for Clk_period;
		Addr <=  "0010010111110";
		Trees_din <= x"ffe2130d";
		wait for Clk_period;
		Addr <=  "0010010111111";
		Trees_din <= x"00db130d";
		wait for Clk_period;
		Addr <=  "0010011000000";
		Trees_din <= x"1800a704";
		wait for Clk_period;
		Addr <=  "0010011000001";
		Trees_din <= x"ff43130d";
		wait for Clk_period;
		Addr <=  "0010011000010";
		Trees_din <= x"0026130d";
		wait for Clk_period;
		Addr <=  "0010011000011";
		Trees_din <= x"03057d44";
		wait for Clk_period;
		Addr <=  "0010011000100";
		Trees_din <= x"040b2b28";
		wait for Clk_period;
		Addr <=  "0010011000101";
		Trees_din <= x"06f2b208";
		wait for Clk_period;
		Addr <=  "0010011000110";
		Trees_din <= x"09003604";
		wait for Clk_period;
		Addr <=  "0010011000111";
		Trees_din <= x"000c13a9";
		wait for Clk_period;
		Addr <=  "0010011001000";
		Trees_din <= x"ff7913a9";
		wait for Clk_period;
		Addr <=  "0010011001001";
		Trees_din <= x"05ff4710";
		wait for Clk_period;
		Addr <=  "0010011001010";
		Trees_din <= x"07ff7108";
		wait for Clk_period;
		Addr <=  "0010011001011";
		Trees_din <= x"05fd6f04";
		wait for Clk_period;
		Addr <=  "0010011001100";
		Trees_din <= x"003813a9";
		wait for Clk_period;
		Addr <=  "0010011001101";
		Trees_din <= x"000113a9";
		wait for Clk_period;
		Addr <=  "0010011001110";
		Trees_din <= x"04048004";
		wait for Clk_period;
		Addr <=  "0010011001111";
		Trees_din <= x"ffd113a9";
		wait for Clk_period;
		Addr <=  "0010011010000";
		Trees_din <= x"000713a9";
		wait for Clk_period;
		Addr <=  "0010011010001";
		Trees_din <= x"14003908";
		wait for Clk_period;
		Addr <=  "0010011010010";
		Trees_din <= x"07010604";
		wait for Clk_period;
		Addr <=  "0010011010011";
		Trees_din <= x"00b013a9";
		wait for Clk_period;
		Addr <=  "0010011010100";
		Trees_din <= x"ff9513a9";
		wait for Clk_period;
		Addr <=  "0010011010101";
		Trees_din <= x"14003f04";
		wait for Clk_period;
		Addr <=  "0010011010110";
		Trees_din <= x"ffaa13a9";
		wait for Clk_period;
		Addr <=  "0010011010111";
		Trees_din <= x"003513a9";
		wait for Clk_period;
		Addr <=  "0010011011000";
		Trees_din <= x"0100630c";
		wait for Clk_period;
		Addr <=  "0010011011001";
		Trees_din <= x"0a022808";
		wait for Clk_period;
		Addr <=  "0010011011010";
		Trees_din <= x"1d023f04";
		wait for Clk_period;
		Addr <=  "0010011011011";
		Trees_din <= x"000713a9";
		wait for Clk_period;
		Addr <=  "0010011011100";
		Trees_din <= x"009113a9";
		wait for Clk_period;
		Addr <=  "0010011011101";
		Trees_din <= x"fff313a9";
		wait for Clk_period;
		Addr <=  "0010011011110";
		Trees_din <= x"040d9708";
		wait for Clk_period;
		Addr <=  "0010011011111";
		Trees_din <= x"1c026f04";
		wait for Clk_period;
		Addr <=  "0010011100000";
		Trees_din <= x"ff9713a9";
		wait for Clk_period;
		Addr <=  "0010011100001";
		Trees_din <= x"002d13a9";
		wait for Clk_period;
		Addr <=  "0010011100010";
		Trees_din <= x"09004804";
		wait for Clk_period;
		Addr <=  "0010011100011";
		Trees_din <= x"008013a9";
		wait for Clk_period;
		Addr <=  "0010011100100";
		Trees_din <= x"fffa13a9";
		wait for Clk_period;
		Addr <=  "0010011100101";
		Trees_din <= x"07f99908";
		wait for Clk_period;
		Addr <=  "0010011100110";
		Trees_din <= x"04fc6604";
		wait for Clk_period;
		Addr <=  "0010011100111";
		Trees_din <= x"ffa413a9";
		wait for Clk_period;
		Addr <=  "0010011101000";
		Trees_din <= x"007213a9";
		wait for Clk_period;
		Addr <=  "0010011101001";
		Trees_din <= x"ff7413a9";
		wait for Clk_period;
		Addr <=  "0010011101010";
		Trees_din <= x"02fd814c";
		wait for Clk_period;
		Addr <=  "0010011101011";
		Trees_din <= x"1f028840";
		wait for Clk_period;
		Addr <=  "0010011101100";
		Trees_din <= x"0c02b620";
		wait for Clk_period;
		Addr <=  "0010011101101";
		Trees_din <= x"12005f10";
		wait for Clk_period;
		Addr <=  "0010011101110";
		Trees_din <= x"13006908";
		wait for Clk_period;
		Addr <=  "0010011101111";
		Trees_din <= x"07fe3904";
		wait for Clk_period;
		Addr <=  "0010011110000";
		Trees_din <= x"ff74149d";
		wait for Clk_period;
		Addr <=  "0010011110001";
		Trees_din <= x"007b149d";
		wait for Clk_period;
		Addr <=  "0010011110010";
		Trees_din <= x"05fb3404";
		wait for Clk_period;
		Addr <=  "0010011110011";
		Trees_din <= x"0066149d";
		wait for Clk_period;
		Addr <=  "0010011110100";
		Trees_din <= x"0006149d";
		wait for Clk_period;
		Addr <=  "0010011110101";
		Trees_din <= x"00ff4708";
		wait for Clk_period;
		Addr <=  "0010011110110";
		Trees_din <= x"03faa504";
		wait for Clk_period;
		Addr <=  "0010011110111";
		Trees_din <= x"fffe149d";
		wait for Clk_period;
		Addr <=  "0010011111000";
		Trees_din <= x"ff4a149d";
		wait for Clk_period;
		Addr <=  "0010011111001";
		Trees_din <= x"02fa1204";
		wait for Clk_period;
		Addr <=  "0010011111010";
		Trees_din <= x"006d149d";
		wait for Clk_period;
		Addr <=  "0010011111011";
		Trees_din <= x"ffbe149d";
		wait for Clk_period;
		Addr <=  "0010011111100";
		Trees_din <= x"00fce810";
		wait for Clk_period;
		Addr <=  "0010011111101";
		Trees_din <= x"05fe2b08";
		wait for Clk_period;
		Addr <=  "0010011111110";
		Trees_din <= x"16034d04";
		wait for Clk_period;
		Addr <=  "0010011111111";
		Trees_din <= x"fffa149d";
		wait for Clk_period;
		Addr <=  "0010100000000";
		Trees_din <= x"ff34149d";
		wait for Clk_period;
		Addr <=  "0010100000001";
		Trees_din <= x"04049404";
		wait for Clk_period;
		Addr <=  "0010100000010";
		Trees_din <= x"ff9b149d";
		wait for Clk_period;
		Addr <=  "0010100000011";
		Trees_din <= x"00d1149d";
		wait for Clk_period;
		Addr <=  "0010100000100";
		Trees_din <= x"10004e08";
		wait for Clk_period;
		Addr <=  "0010100000101";
		Trees_din <= x"11000204";
		wait for Clk_period;
		Addr <=  "0010100000110";
		Trees_din <= x"0049149d";
		wait for Clk_period;
		Addr <=  "0010100000111";
		Trees_din <= x"ff54149d";
		wait for Clk_period;
		Addr <=  "0010100001000";
		Trees_din <= x"0b00eb04";
		wait for Clk_period;
		Addr <=  "0010100001001";
		Trees_din <= x"006b149d";
		wait for Clk_period;
		Addr <=  "0010100001010";
		Trees_din <= x"ff96149d";
		wait for Clk_period;
		Addr <=  "0010100001011";
		Trees_din <= x"00fce804";
		wait for Clk_period;
		Addr <=  "0010100001100";
		Trees_din <= x"0071149d";
		wait for Clk_period;
		Addr <=  "0010100001101";
		Trees_din <= x"1002b304";
		wait for Clk_period;
		Addr <=  "0010100001110";
		Trees_din <= x"ff33149d";
		wait for Clk_period;
		Addr <=  "0010100001111";
		Trees_din <= x"002b149d";
		wait for Clk_period;
		Addr <=  "0010100010000";
		Trees_din <= x"0e004128";
		wait for Clk_period;
		Addr <=  "0010100010001";
		Trees_din <= x"0d006610";
		wait for Clk_period;
		Addr <=  "0010100010010";
		Trees_din <= x"0c01cd0c";
		wait for Clk_period;
		Addr <=  "0010100010011";
		Trees_din <= x"15f73e04";
		wait for Clk_period;
		Addr <=  "0010100010100";
		Trees_din <= x"fff0149d";
		wait for Clk_period;
		Addr <=  "0010100010101";
		Trees_din <= x"0c013c04";
		wait for Clk_period;
		Addr <=  "0010100010110";
		Trees_din <= x"0124149d";
		wait for Clk_period;
		Addr <=  "0010100010111";
		Trees_din <= x"0045149d";
		wait for Clk_period;
		Addr <=  "0010100011000";
		Trees_din <= x"ffef149d";
		wait for Clk_period;
		Addr <=  "0010100011001";
		Trees_din <= x"1f024d0c";
		wait for Clk_period;
		Addr <=  "0010100011010";
		Trees_din <= x"0b00b404";
		wait for Clk_period;
		Addr <=  "0010100011011";
		Trees_din <= x"0008149d";
		wait for Clk_period;
		Addr <=  "0010100011100";
		Trees_din <= x"02ff5e04";
		wait for Clk_period;
		Addr <=  "0010100011101";
		Trees_din <= x"ff34149d";
		wait for Clk_period;
		Addr <=  "0010100011110";
		Trees_din <= x"ffc1149d";
		wait for Clk_period;
		Addr <=  "0010100011111";
		Trees_din <= x"18005404";
		wait for Clk_period;
		Addr <=  "0010100100000";
		Trees_din <= x"ff71149d";
		wait for Clk_period;
		Addr <=  "0010100100001";
		Trees_din <= x"02fda804";
		wait for Clk_period;
		Addr <=  "0010100100010";
		Trees_din <= x"ff85149d";
		wait for Clk_period;
		Addr <=  "0010100100011";
		Trees_din <= x"001e149d";
		wait for Clk_period;
		Addr <=  "0010100100100";
		Trees_din <= x"1800a704";
		wait for Clk_period;
		Addr <=  "0010100100101";
		Trees_din <= x"ff4c149d";
		wait for Clk_period;
		Addr <=  "0010100100110";
		Trees_din <= x"0021149d";
		wait for Clk_period;
		Addr <=  "0010100100111";
		Trees_din <= x"04fb9604";
		wait for Clk_period;
		Addr <=  "0010100101000";
		Trees_din <= x"ff831531";
		wait for Clk_period;
		Addr <=  "0010100101001";
		Trees_din <= x"21000128";
		wait for Clk_period;
		Addr <=  "0010100101010";
		Trees_din <= x"21000120";
		wait for Clk_period;
		Addr <=  "0010100101011";
		Trees_din <= x"040ab810";
		wait for Clk_period;
		Addr <=  "0010100101100";
		Trees_din <= x"01fd9608";
		wait for Clk_period;
		Addr <=  "0010100101101";
		Trees_din <= x"060c0004";
		wait for Clk_period;
		Addr <=  "0010100101110";
		Trees_din <= x"00161531";
		wait for Clk_period;
		Addr <=  "0010100101111";
		Trees_din <= x"ff8a1531";
		wait for Clk_period;
		Addr <=  "0010100110000";
		Trees_din <= x"060b8504";
		wait for Clk_period;
		Addr <=  "0010100110001";
		Trees_din <= x"fffa1531";
		wait for Clk_period;
		Addr <=  "0010100110010";
		Trees_din <= x"004f1531";
		wait for Clk_period;
		Addr <=  "0010100110011";
		Trees_din <= x"0e004a08";
		wait for Clk_period;
		Addr <=  "0010100110100";
		Trees_din <= x"15f76804";
		wait for Clk_period;
		Addr <=  "0010100110101";
		Trees_din <= x"00001531";
		wait for Clk_period;
		Addr <=  "0010100110110";
		Trees_din <= x"006c1531";
		wait for Clk_period;
		Addr <=  "0010100110111";
		Trees_din <= x"03fb5a04";
		wait for Clk_period;
		Addr <=  "0010100111000";
		Trees_din <= x"00251531";
		wait for Clk_period;
		Addr <=  "0010100111001";
		Trees_din <= x"ff971531";
		wait for Clk_period;
		Addr <=  "0010100111010";
		Trees_din <= x"00fed004";
		wait for Clk_period;
		Addr <=  "0010100111011";
		Trees_din <= x"00fb1531";
		wait for Clk_period;
		Addr <=  "0010100111100";
		Trees_din <= x"002a1531";
		wait for Clk_period;
		Addr <=  "0010100111101";
		Trees_din <= x"18005008";
		wait for Clk_period;
		Addr <=  "0010100111110";
		Trees_din <= x"01fe2904";
		wait for Clk_period;
		Addr <=  "0010100111111";
		Trees_din <= x"ffbf1531";
		wait for Clk_period;
		Addr <=  "0010101000000";
		Trees_din <= x"00b31531";
		wait for Clk_period;
		Addr <=  "0010101000001";
		Trees_din <= x"0d006f08";
		wait for Clk_period;
		Addr <=  "0010101000010";
		Trees_din <= x"0d006d04";
		wait for Clk_period;
		Addr <=  "0010101000011";
		Trees_din <= x"00001531";
		wait for Clk_period;
		Addr <=  "0010101000100";
		Trees_din <= x"00981531";
		wait for Clk_period;
		Addr <=  "0010101000101";
		Trees_din <= x"0b006008";
		wait for Clk_period;
		Addr <=  "0010101000110";
		Trees_din <= x"04050004";
		wait for Clk_period;
		Addr <=  "0010101000111";
		Trees_din <= x"ff911531";
		wait for Clk_period;
		Addr <=  "0010101001000";
		Trees_din <= x"004c1531";
		wait for Clk_period;
		Addr <=  "0010101001001";
		Trees_din <= x"06050904";
		wait for Clk_period;
		Addr <=  "0010101001010";
		Trees_din <= x"ffd01531";
		wait for Clk_period;
		Addr <=  "0010101001011";
		Trees_din <= x"ff451531";
		wait for Clk_period;
		Addr <=  "0010101001100";
		Trees_din <= x"03057d58";
		wait for Clk_period;
		Addr <=  "0010101001101";
		Trees_din <= x"0b004b28";
		wait for Clk_period;
		Addr <=  "0010101001110";
		Trees_din <= x"08005218";
		wait for Clk_period;
		Addr <=  "0010101001111";
		Trees_din <= x"0a02eb10";
		wait for Clk_period;
		Addr <=  "0010101010000";
		Trees_din <= x"1100b808";
		wait for Clk_period;
		Addr <=  "0010101010001";
		Trees_din <= x"00fdd604";
		wait for Clk_period;
		Addr <=  "0010101010010";
		Trees_din <= x"006615f5";
		wait for Clk_period;
		Addr <=  "0010101010011";
		Trees_din <= x"fff215f5";
		wait for Clk_period;
		Addr <=  "0010101010100";
		Trees_din <= x"1e028704";
		wait for Clk_period;
		Addr <=  "0010101010101";
		Trees_din <= x"00ea15f5";
		wait for Clk_period;
		Addr <=  "0010101010110";
		Trees_din <= x"003815f5";
		wait for Clk_period;
		Addr <=  "0010101010111";
		Trees_din <= x"17011f04";
		wait for Clk_period;
		Addr <=  "0010101011000";
		Trees_din <= x"006b15f5";
		wait for Clk_period;
		Addr <=  "0010101011001";
		Trees_din <= x"ff9b15f5";
		wait for Clk_period;
		Addr <=  "0010101011010";
		Trees_din <= x"1c028308";
		wait for Clk_period;
		Addr <=  "0010101011011";
		Trees_din <= x"0d009f04";
		wait for Clk_period;
		Addr <=  "0010101011100";
		Trees_din <= x"ffcb15f5";
		wait for Clk_period;
		Addr <=  "0010101011101";
		Trees_din <= x"00ab15f5";
		wait for Clk_period;
		Addr <=  "0010101011110";
		Trees_din <= x"06072d04";
		wait for Clk_period;
		Addr <=  "0010101011111";
		Trees_din <= x"002515f5";
		wait for Clk_period;
		Addr <=  "0010101100000";
		Trees_din <= x"ff5715f5";
		wait for Clk_period;
		Addr <=  "0010101100001";
		Trees_din <= x"08003810";
		wait for Clk_period;
		Addr <=  "0010101100010";
		Trees_din <= x"04069a0c";
		wait for Clk_period;
		Addr <=  "0010101100011";
		Trees_din <= x"0d004e08";
		wait for Clk_period;
		Addr <=  "0010101100100";
		Trees_din <= x"0a000204";
		wait for Clk_period;
		Addr <=  "0010101100101";
		Trees_din <= x"ff9f15f5";
		wait for Clk_period;
		Addr <=  "0010101100110";
		Trees_din <= x"006f15f5";
		wait for Clk_period;
		Addr <=  "0010101100111";
		Trees_din <= x"ff5615f5";
		wait for Clk_period;
		Addr <=  "0010101101000";
		Trees_din <= x"007d15f5";
		wait for Clk_period;
		Addr <=  "0010101101001";
		Trees_din <= x"21000110";
		wait for Clk_period;
		Addr <=  "0010101101010";
		Trees_din <= x"21000108";
		wait for Clk_period;
		Addr <=  "0010101101011";
		Trees_din <= x"08003b04";
		wait for Clk_period;
		Addr <=  "0010101101100";
		Trees_din <= x"004015f5";
		wait for Clk_period;
		Addr <=  "0010101101101";
		Trees_din <= x"000615f5";
		wait for Clk_period;
		Addr <=  "0010101101110";
		Trees_din <= x"00fed004";
		wait for Clk_period;
		Addr <=  "0010101101111";
		Trees_din <= x"00e315f5";
		wait for Clk_period;
		Addr <=  "0010101110000";
		Trees_din <= x"002715f5";
		wait for Clk_period;
		Addr <=  "0010101110001";
		Trees_din <= x"0d006f08";
		wait for Clk_period;
		Addr <=  "0010101110010";
		Trees_din <= x"0d006d04";
		wait for Clk_period;
		Addr <=  "0010101110011";
		Trees_din <= x"000015f5";
		wait for Clk_period;
		Addr <=  "0010101110100";
		Trees_din <= x"009115f5";
		wait for Clk_period;
		Addr <=  "0010101110101";
		Trees_din <= x"18005004";
		wait for Clk_period;
		Addr <=  "0010101110110";
		Trees_din <= x"005615f5";
		wait for Clk_period;
		Addr <=  "0010101110111";
		Trees_din <= x"ff6f15f5";
		wait for Clk_period;
		Addr <=  "0010101111000";
		Trees_din <= x"07f99908";
		wait for Clk_period;
		Addr <=  "0010101111001";
		Trees_din <= x"06029204";
		wait for Clk_period;
		Addr <=  "0010101111010";
		Trees_din <= x"ffec15f5";
		wait for Clk_period;
		Addr <=  "0010101111011";
		Trees_din <= x"003a15f5";
		wait for Clk_period;
		Addr <=  "0010101111100";
		Trees_din <= x"ff7915f5";
		wait for Clk_period;
		Addr <=  "0010101111101";
		Trees_din <= x"02fd8148";
		wait for Clk_period;
		Addr <=  "0010101111110";
		Trees_din <= x"1f02883c";
		wait for Clk_period;
		Addr <=  "0010101111111";
		Trees_din <= x"07fedb1c";
		wait for Clk_period;
		Addr <=  "0010110000000";
		Trees_din <= x"02f9c10c";
		wait for Clk_period;
		Addr <=  "0010110000001";
		Trees_din <= x"04047904";
		wait for Clk_period;
		Addr <=  "0010110000010";
		Trees_din <= x"ffac16e1";
		wait for Clk_period;
		Addr <=  "0010110000011";
		Trees_din <= x"05fd9104";
		wait for Clk_period;
		Addr <=  "0010110000100";
		Trees_din <= x"00eb16e1";
		wait for Clk_period;
		Addr <=  "0010110000101";
		Trees_din <= x"001816e1";
		wait for Clk_period;
		Addr <=  "0010110000110";
		Trees_din <= x"09004208";
		wait for Clk_period;
		Addr <=  "0010110000111";
		Trees_din <= x"09003504";
		wait for Clk_period;
		Addr <=  "0010110001000";
		Trees_din <= x"ffe216e1";
		wait for Clk_period;
		Addr <=  "0010110001001";
		Trees_din <= x"004a16e1";
		wait for Clk_period;
		Addr <=  "0010110001010";
		Trees_din <= x"05fd6f04";
		wait for Clk_period;
		Addr <=  "0010110001011";
		Trees_din <= x"003f16e1";
		wait for Clk_period;
		Addr <=  "0010110001100";
		Trees_din <= x"ffc116e1";
		wait for Clk_period;
		Addr <=  "0010110001101";
		Trees_din <= x"1f028510";
		wait for Clk_period;
		Addr <=  "0010110001110";
		Trees_din <= x"0f008008";
		wait for Clk_period;
		Addr <=  "0010110001111";
		Trees_din <= x"0408c104";
		wait for Clk_period;
		Addr <=  "0010110010000";
		Trees_din <= x"000216e1";
		wait for Clk_period;
		Addr <=  "0010110010001";
		Trees_din <= x"004016e1";
		wait for Clk_period;
		Addr <=  "0010110010010";
		Trees_din <= x"0b00a004";
		wait for Clk_period;
		Addr <=  "0010110010011";
		Trees_din <= x"000b16e1";
		wait for Clk_period;
		Addr <=  "0010110010100";
		Trees_din <= x"ffba16e1";
		wait for Clk_period;
		Addr <=  "0010110010101";
		Trees_din <= x"0a000b08";
		wait for Clk_period;
		Addr <=  "0010110010110";
		Trees_din <= x"02fb1604";
		wait for Clk_period;
		Addr <=  "0010110010111";
		Trees_din <= x"ff5216e1";
		wait for Clk_period;
		Addr <=  "0010110011000";
		Trees_din <= x"007d16e1";
		wait for Clk_period;
		Addr <=  "0010110011001";
		Trees_din <= x"18005f04";
		wait for Clk_period;
		Addr <=  "0010110011010";
		Trees_din <= x"00af16e1";
		wait for Clk_period;
		Addr <=  "0010110011011";
		Trees_din <= x"000d16e1";
		wait for Clk_period;
		Addr <=  "0010110011100";
		Trees_din <= x"00fce804";
		wait for Clk_period;
		Addr <=  "0010110011101";
		Trees_din <= x"006916e1";
		wait for Clk_period;
		Addr <=  "0010110011110";
		Trees_din <= x"1002b304";
		wait for Clk_period;
		Addr <=  "0010110011111";
		Trees_din <= x"ff3f16e1";
		wait for Clk_period;
		Addr <=  "0010110100000";
		Trees_din <= x"002b16e1";
		wait for Clk_period;
		Addr <=  "0010110100001";
		Trees_din <= x"0e004128";
		wait for Clk_period;
		Addr <=  "0010110100010";
		Trees_din <= x"0d006610";
		wait for Clk_period;
		Addr <=  "0010110100011";
		Trees_din <= x"0f006e08";
		wait for Clk_period;
		Addr <=  "0010110100100";
		Trees_din <= x"02fe9304";
		wait for Clk_period;
		Addr <=  "0010110100101";
		Trees_din <= x"00f316e1";
		wait for Clk_period;
		Addr <=  "0010110100110";
		Trees_din <= x"fffe16e1";
		wait for Clk_period;
		Addr <=  "0010110100111";
		Trees_din <= x"11011d04";
		wait for Clk_period;
		Addr <=  "0010110101000";
		Trees_din <= x"ffc016e1";
		wait for Clk_period;
		Addr <=  "0010110101001";
		Trees_din <= x"005716e1";
		wait for Clk_period;
		Addr <=  "0010110101010";
		Trees_din <= x"0b00ef10";
		wait for Clk_period;
		Addr <=  "0010110101011";
		Trees_din <= x"0b00e808";
		wait for Clk_period;
		Addr <=  "0010110101100";
		Trees_din <= x"07004104";
		wait for Clk_period;
		Addr <=  "0010110101101";
		Trees_din <= x"ffca16e1";
		wait for Clk_period;
		Addr <=  "0010110101110";
		Trees_din <= x"003a16e1";
		wait for Clk_period;
		Addr <=  "0010110101111";
		Trees_din <= x"0a006d04";
		wait for Clk_period;
		Addr <=  "0010110110000";
		Trees_din <= x"000116e1";
		wait for Clk_period;
		Addr <=  "0010110110001";
		Trees_din <= x"010616e1";
		wait for Clk_period;
		Addr <=  "0010110110010";
		Trees_din <= x"18005d04";
		wait for Clk_period;
		Addr <=  "0010110110011";
		Trees_din <= x"001a16e1";
		wait for Clk_period;
		Addr <=  "0010110110100";
		Trees_din <= x"ff3416e1";
		wait for Clk_period;
		Addr <=  "0010110110101";
		Trees_din <= x"08004d04";
		wait for Clk_period;
		Addr <=  "0010110110110";
		Trees_din <= x"ff5316e1";
		wait for Clk_period;
		Addr <=  "0010110110111";
		Trees_din <= x"fff816e1";
		wait for Clk_period;
		Addr <=  "0010110111000";
		Trees_din <= x"03057d78";
		wait for Clk_period;
		Addr <=  "0010110111001";
		Trees_din <= x"0d00883c";
		wait for Clk_period;
		Addr <=  "0010110111010";
		Trees_din <= x"08004f20";
		wait for Clk_period;
		Addr <=  "0010110111011";
		Trees_din <= x"0b009710";
		wait for Clk_period;
		Addr <=  "0010110111100";
		Trees_din <= x"0404d308";
		wait for Clk_period;
		Addr <=  "0010110111101";
		Trees_din <= x"03fece04";
		wait for Clk_period;
		Addr <=  "0010110111110";
		Trees_din <= x"ff7617e5";
		wait for Clk_period;
		Addr <=  "0010110111111";
		Trees_din <= x"003917e5";
		wait for Clk_period;
		Addr <=  "0010111000000";
		Trees_din <= x"0f008804";
		wait for Clk_period;
		Addr <=  "0010111000001";
		Trees_din <= x"008917e5";
		wait for Clk_period;
		Addr <=  "0010111000010";
		Trees_din <= x"ffba17e5";
		wait for Clk_period;
		Addr <=  "0010111000011";
		Trees_din <= x"0b009d08";
		wait for Clk_period;
		Addr <=  "0010111000100";
		Trees_din <= x"04082404";
		wait for Clk_period;
		Addr <=  "0010111000101";
		Trees_din <= x"ff8117e5";
		wait for Clk_period;
		Addr <=  "0010111000110";
		Trees_din <= x"007017e5";
		wait for Clk_period;
		Addr <=  "0010111000111";
		Trees_din <= x"12005304";
		wait for Clk_period;
		Addr <=  "0010111001000";
		Trees_din <= x"000017e5";
		wait for Clk_period;
		Addr <=  "0010111001001";
		Trees_din <= x"004917e5";
		wait for Clk_period;
		Addr <=  "0010111001010";
		Trees_din <= x"0f008810";
		wait for Clk_period;
		Addr <=  "0010111001011";
		Trees_din <= x"1300af08";
		wait for Clk_period;
		Addr <=  "0010111001100";
		Trees_din <= x"05fe1f04";
		wait for Clk_period;
		Addr <=  "0010111001101";
		Trees_din <= x"ffb917e5";
		wait for Clk_period;
		Addr <=  "0010111001110";
		Trees_din <= x"002517e5";
		wait for Clk_period;
		Addr <=  "0010111001111";
		Trees_din <= x"07fd6a04";
		wait for Clk_period;
		Addr <=  "0010111010000";
		Trees_din <= x"001a17e5";
		wait for Clk_period;
		Addr <=  "0010111010001";
		Trees_din <= x"ff0717e5";
		wait for Clk_period;
		Addr <=  "0010111010010";
		Trees_din <= x"00fea408";
		wait for Clk_period;
		Addr <=  "0010111010011";
		Trees_din <= x"0c014604";
		wait for Clk_period;
		Addr <=  "0010111010100";
		Trees_din <= x"004517e5";
		wait for Clk_period;
		Addr <=  "0010111010101";
		Trees_din <= x"ff7c17e5";
		wait for Clk_period;
		Addr <=  "0010111010110";
		Trees_din <= x"00e217e5";
		wait for Clk_period;
		Addr <=  "0010111010111";
		Trees_din <= x"00fd1520";
		wait for Clk_period;
		Addr <=  "0010111011000";
		Trees_din <= x"00fc7f10";
		wait for Clk_period;
		Addr <=  "0010111011001";
		Trees_din <= x"1b027408";
		wait for Clk_period;
		Addr <=  "0010111011010";
		Trees_din <= x"1f024004";
		wait for Clk_period;
		Addr <=  "0010111011011";
		Trees_din <= x"007c17e5";
		wait for Clk_period;
		Addr <=  "0010111011100";
		Trees_din <= x"000f17e5";
		wait for Clk_period;
		Addr <=  "0010111011101";
		Trees_din <= x"11006204";
		wait for Clk_period;
		Addr <=  "0010111011110";
		Trees_din <= x"ff6317e5";
		wait for Clk_period;
		Addr <=  "0010111011111";
		Trees_din <= x"ffeb17e5";
		wait for Clk_period;
		Addr <=  "0010111100000";
		Trees_din <= x"01fe8808";
		wait for Clk_period;
		Addr <=  "0010111100001";
		Trees_din <= x"1703de04";
		wait for Clk_period;
		Addr <=  "0010111100010";
		Trees_din <= x"010017e5";
		wait for Clk_period;
		Addr <=  "0010111100011";
		Trees_din <= x"003817e5";
		wait for Clk_period;
		Addr <=  "0010111100100";
		Trees_din <= x"0604e204";
		wait for Clk_period;
		Addr <=  "0010111100101";
		Trees_din <= x"007917e5";
		wait for Clk_period;
		Addr <=  "0010111100110";
		Trees_din <= x"ffa817e5";
		wait for Clk_period;
		Addr <=  "0010111100111";
		Trees_din <= x"00feff0c";
		wait for Clk_period;
		Addr <=  "0010111101000";
		Trees_din <= x"0a03e708";
		wait for Clk_period;
		Addr <=  "0010111101001";
		Trees_din <= x"0609be04";
		wait for Clk_period;
		Addr <=  "0010111101010";
		Trees_din <= x"000717e5";
		wait for Clk_period;
		Addr <=  "0010111101011";
		Trees_din <= x"ffa817e5";
		wait for Clk_period;
		Addr <=  "0010111101100";
		Trees_din <= x"00d917e5";
		wait for Clk_period;
		Addr <=  "0010111101101";
		Trees_din <= x"03fcf908";
		wait for Clk_period;
		Addr <=  "0010111101110";
		Trees_din <= x"07006004";
		wait for Clk_period;
		Addr <=  "0010111101111";
		Trees_din <= x"010317e5";
		wait for Clk_period;
		Addr <=  "0010111110000";
		Trees_din <= x"004017e5";
		wait for Clk_period;
		Addr <=  "0010111110001";
		Trees_din <= x"09002e04";
		wait for Clk_period;
		Addr <=  "0010111110010";
		Trees_din <= x"009617e5";
		wait for Clk_period;
		Addr <=  "0010111110011";
		Trees_din <= x"ffab17e5";
		wait for Clk_period;
		Addr <=  "0010111110100";
		Trees_din <= x"07f99908";
		wait for Clk_period;
		Addr <=  "0010111110101";
		Trees_din <= x"11000c04";
		wait for Clk_period;
		Addr <=  "0010111110110";
		Trees_din <= x"fff317e5";
		wait for Clk_period;
		Addr <=  "0010111110111";
		Trees_din <= x"002b17e5";
		wait for Clk_period;
		Addr <=  "0010111111000";
		Trees_din <= x"ff7d17e5";
		wait for Clk_period;
		Addr <=  "0010111111001";
		Trees_din <= x"05fb341c";
		wait for Clk_period;
		Addr <=  "0010111111010";
		Trees_din <= x"0b00bc0c";
		wait for Clk_period;
		Addr <=  "0010111111011";
		Trees_din <= x"03fb1704";
		wait for Clk_period;
		Addr <=  "0010111111100";
		Trees_din <= x"007518e1";
		wait for Clk_period;
		Addr <=  "0010111111101";
		Trees_din <= x"11000704";
		wait for Clk_period;
		Addr <=  "0010111111110";
		Trees_din <= x"ff5318e1";
		wait for Clk_period;
		Addr <=  "0010111111111";
		Trees_din <= x"fff618e1";
		wait for Clk_period;
		Addr <=  "0011000000000";
		Trees_din <= x"07000e04";
		wait for Clk_period;
		Addr <=  "0011000000001";
		Trees_din <= x"ffdc18e1";
		wait for Clk_period;
		Addr <=  "0011000000010";
		Trees_din <= x"1300b508";
		wait for Clk_period;
		Addr <=  "0011000000011";
		Trees_din <= x"06fb6604";
		wait for Clk_period;
		Addr <=  "0011000000100";
		Trees_din <= x"003c18e1";
		wait for Clk_period;
		Addr <=  "0011000000101";
		Trees_din <= x"00d418e1";
		wait for Clk_period;
		Addr <=  "0011000000110";
		Trees_din <= x"001b18e1";
		wait for Clk_period;
		Addr <=  "0011000000111";
		Trees_din <= x"03fa3e24";
		wait for Clk_period;
		Addr <=  "0011000001000";
		Trees_din <= x"1afc9e18";
		wait for Clk_period;
		Addr <=  "0011000001001";
		Trees_din <= x"1603f70c";
		wait for Clk_period;
		Addr <=  "0011000001010";
		Trees_din <= x"14004108";
		wait for Clk_period;
		Addr <=  "0011000001011";
		Trees_din <= x"00fd6504";
		wait for Clk_period;
		Addr <=  "0011000001100";
		Trees_din <= x"ff8f18e1";
		wait for Clk_period;
		Addr <=  "0011000001101";
		Trees_din <= x"004b18e1";
		wait for Clk_period;
		Addr <=  "0011000001110";
		Trees_din <= x"ff3518e1";
		wait for Clk_period;
		Addr <=  "0011000001111";
		Trees_din <= x"18006304";
		wait for Clk_period;
		Addr <=  "0011000010000";
		Trees_din <= x"002f18e1";
		wait for Clk_period;
		Addr <=  "0011000010001";
		Trees_din <= x"05fc7304";
		wait for Clk_period;
		Addr <=  "0011000010010";
		Trees_din <= x"003918e1";
		wait for Clk_period;
		Addr <=  "0011000010011";
		Trees_din <= x"00cf18e1";
		wait for Clk_period;
		Addr <=  "0011000010100";
		Trees_din <= x"0a00c808";
		wait for Clk_period;
		Addr <=  "0011000010101";
		Trees_din <= x"15f6e704";
		wait for Clk_period;
		Addr <=  "0011000010110";
		Trees_din <= x"ffec18e1";
		wait for Clk_period;
		Addr <=  "0011000010111";
		Trees_din <= x"ff3f18e1";
		wait for Clk_period;
		Addr <=  "0011000011000";
		Trees_din <= x"002b18e1";
		wait for Clk_period;
		Addr <=  "0011000011001";
		Trees_din <= x"03fabd20";
		wait for Clk_period;
		Addr <=  "0011000011010";
		Trees_din <= x"1e025710";
		wait for Clk_period;
		Addr <=  "0011000011011";
		Trees_din <= x"00fea108";
		wait for Clk_period;
		Addr <=  "0011000011100";
		Trees_din <= x"00fd5304";
		wait for Clk_period;
		Addr <=  "0011000011101";
		Trees_din <= x"005418e1";
		wait for Clk_period;
		Addr <=  "0011000011110";
		Trees_din <= x"00f818e1";
		wait for Clk_period;
		Addr <=  "0011000011111";
		Trees_din <= x"06066c04";
		wait for Clk_period;
		Addr <=  "0011000100000";
		Trees_din <= x"009818e1";
		wait for Clk_period;
		Addr <=  "0011000100001";
		Trees_din <= x"ff6818e1";
		wait for Clk_period;
		Addr <=  "0011000100010";
		Trees_din <= x"02faf208";
		wait for Clk_period;
		Addr <=  "0011000100011";
		Trees_din <= x"07031004";
		wait for Clk_period;
		Addr <=  "0011000100100";
		Trees_din <= x"005218e1";
		wait for Clk_period;
		Addr <=  "0011000100101";
		Trees_din <= x"ffa018e1";
		wait for Clk_period;
		Addr <=  "0011000100110";
		Trees_din <= x"0a00e904";
		wait for Clk_period;
		Addr <=  "0011000100111";
		Trees_din <= x"ffda18e1";
		wait for Clk_period;
		Addr <=  "0011000101000";
		Trees_din <= x"ff4918e1";
		wait for Clk_period;
		Addr <=  "0011000101001";
		Trees_din <= x"1703fa10";
		wait for Clk_period;
		Addr <=  "0011000101010";
		Trees_din <= x"0c006f08";
		wait for Clk_period;
		Addr <=  "0011000101011";
		Trees_din <= x"0b00cb04";
		wait for Clk_period;
		Addr <=  "0011000101100";
		Trees_din <= x"001a18e1";
		wait for Clk_period;
		Addr <=  "0011000101101";
		Trees_din <= x"010118e1";
		wait for Clk_period;
		Addr <=  "0011000101110";
		Trees_din <= x"15f6f004";
		wait for Clk_period;
		Addr <=  "0011000101111";
		Trees_din <= x"008518e1";
		wait for Clk_period;
		Addr <=  "0011000110000";
		Trees_din <= x"000318e1";
		wait for Clk_period;
		Addr <=  "0011000110001";
		Trees_din <= x"0700ca08";
		wait for Clk_period;
		Addr <=  "0011000110010";
		Trees_din <= x"03fcbb04";
		wait for Clk_period;
		Addr <=  "0011000110011";
		Trees_din <= x"003518e1";
		wait for Clk_period;
		Addr <=  "0011000110100";
		Trees_din <= x"ffe518e1";
		wait for Clk_period;
		Addr <=  "0011000110101";
		Trees_din <= x"04069004";
		wait for Clk_period;
		Addr <=  "0011000110110";
		Trees_din <= x"ff9218e1";
		wait for Clk_period;
		Addr <=  "0011000110111";
		Trees_din <= x"fff318e1";
		wait for Clk_period;
		Addr <=  "0011000111000";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  2
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"0304e150";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"03028a1c";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"03ff4708";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"00facd04";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"0000014d";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"ff52014d";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"1bf9f804";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"0070014d";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"05fe1b08";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"03ff6304";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"006d014d";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"ff8a014d";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"08005b04";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"ff5c014d";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"000f014d";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"05ff841c";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"0e00230c";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"1c028508";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"1e026904";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"0070014d";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"029d014d";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"ffa4014d";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"12004d08";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"07fe3004";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"ff77014d";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"006b014d";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"05fe5704";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"018d014d";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"ffd6014d";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"07ff980c";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"09002004";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"0037014d";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"09004b04";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"ff56014d";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"000f014d";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"04fae404";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"ff79014d";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"08004804";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"015c014d";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"ff9c014d";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"05020f34";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"0307f81c";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"060ada0c";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"0207e908";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"16040004";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"0282014d";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"ffa4014d";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"ff9c014d";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"03067c08";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"09003404";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"00ca014d";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"ff8a014d";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"05ffa104";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"ffce014d";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"026e014d";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"060ada08";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"01004704";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"0462014d";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"0037014d";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"01fcbc08";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"08004904";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"ff90014d";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"00ca014d";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"0309a404";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"00a6014d";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"0304014d";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"06f9a108";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"00fc7f04";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"0021014d";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"ff54014d";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"030c5010";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"04fb4b08";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"01fbc904";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"00a6014d";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"ff7e014d";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"060ac504";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"0282014d";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"0037014d";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"04e87804";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"ff84014d";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"1100ae04";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"03ae014d";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"00ca014d";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"03030730";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"03ff4708";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"00facd04";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"00090239";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"ff570239";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"1e02871c";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"08003c0c";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"05fe5108";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"08003b04";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"ff810239";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"01210239";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"ff6f0239";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"0a001508";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"12004404";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"00050239";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"ff780239";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"0c032f04";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"ff600239";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"ffc30239";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"17029204";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"01500239";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"03028a04";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"ff700239";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"00be0239";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"05063430";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"03067c1c";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"07fdfa10";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"0d007908";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"0f005a04";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"00610239";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"ff6a0239";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"1300b904";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"01360239";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"ffe30239";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"08003e04";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"ff790239";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"06097f04";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"016d0239";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"00230239";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"0209ce10";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"060d4208";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"0001e004";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"01c10239";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"00450239";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"0309a404";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"ff700239";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"013a0239";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"ff790239";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"06f53804";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"ff5b0239";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"03093c08";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"0f008c04";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"ff610239";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"00110239";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"05157908";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"0609ff04";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"018a0239";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"ffa80239";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"ff770239";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"03030734";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"03ff4708";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"00facd04";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"000f031d";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"ff5b031d";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"1e02871c";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"03ff630c";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"06068d08";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"15f73904";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"015c031d";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"001c031d";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"ff75031d";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"08003c08";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"0c026a04";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"ffac031d";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"00b6031d";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"09003304";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"ffc5031d";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"ff6e031d";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"09003d04";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"ff7e031d";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"05ff4d08";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"02fc2b04";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"0023031d";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"0189031d";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"ff9c031d";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"05063424";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"03067c10";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"1d02840c";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"02021c08";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"060ada04";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"00d9031d";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"ffef031d";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"ff6d031d";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"ff65031d";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"0209ce10";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"060d4208";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"18003f04";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"0018031d";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"012f031d";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"0309a404";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"ff78031d";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"00df031d";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"ff82031d";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"06f53804";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"ff5f031d";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"08004310";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"0308dd08";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"19000604";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"ff80031d";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"0041031d";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"04e87804";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"ff9b031d";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"015d031d";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"10000104";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"0003031d";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"ff66031d";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"03030738";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"03ff4708";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"00facd04";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"00150409";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"ff5e0409";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"1e028720";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"0a002710";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"12004408";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"05ff0804";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"00890409";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"ff700409";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"05fc8004";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"00920409";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"ff760409";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"08003c08";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"11001504";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"00bf0409";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"ffa00409";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"0c032f04";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"ff660409";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"ffe40409";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"14003a04";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"ff850409";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"0a004104";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"ff9c0409";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"0300cf04";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"000a0409";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"01760409";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"0101b430";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"0305fb18";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"04fe810c";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"18007104";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"ff620409";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"01fcdf04";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"00e70409";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"ffbd0409";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"1d028408";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"1f026404";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"001a0409";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"00fe0409";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"ff760409";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"02fef00c";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"06105808";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"14004f04";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"00f60409";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"fffa0409";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"ff9c0409";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"060d3208";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"09004704";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"00a70409";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"ffa10409";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"ff730409";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"06f9a104";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"ff620409";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"0a001708";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"15f74704";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"00040409";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"00ac0409";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"ff840409";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"03028a3c";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"03ff4710";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"00facd04";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"001a0505";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"11033504";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"ff5f0505";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"0e004604";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"ff770505";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"00470505";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"04020c10";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"0c02d808";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"2003ff04";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"fff70505";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"ff600505";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"12004204";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"00d80505";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"ff810505";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"1f02430c";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"0f007104";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"ff8e0505";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"11018204";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"01800505";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"ffa10505";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"0a000708";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"0b00d604";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"ff7d0505";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"00f90505";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"01fc8604";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"00320505";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"ff7c0505";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"0506342c";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"0307f81c";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"060d4210";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"02021c08";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"0d007904";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"002a0505";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"00a60505";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"15f6f504";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"00140505";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"ff710505";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"01fba504";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"00ca0505";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"18009404";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"ff680505";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"00450505";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"0209ce0c";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"1d028808";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"0e004904";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"00cf0505";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"fff10505";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"ffd30505";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"ff9f0505";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"06f53804";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"ff660505";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"03093c08";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"19001704";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"ff6a0505";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"002f0505";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"0f007708";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"04e87804";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"ffaa0505";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"00f30505";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"ff890505";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"03028a3c";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"03ff4710";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"00facd04";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"001f0611";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"11033504";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"ff610611";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"15fa7f04";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"00480611";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"ff7b0611";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"04020c10";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"0c02d808";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"2003ff04";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"fffc0611";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"ff630611";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"12004204";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"00bb0611";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"ff870611";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"12004510";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"11000608";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"0d008204";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"016c0611";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"ffa10611";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"01fd2504";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"00aa0611";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"ffb00611";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"04022f04";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"00bd0611";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"14004d04";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"ff640611";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"000d0611";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"01020b40";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"0305fb20";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"05006210";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"08004108";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"1afc0104";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"004b0611";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"ff7f0611";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"02fc4e04";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"000d0611";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"00bd0611";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"0e003908";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"02fbab04";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"001f0611";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"ff640611";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"07fd6a04";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"ff830611";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"007c0611";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"02fef010";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"0d007a08";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"060ac504";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"00a80611";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"00180611";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"1a013e04";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"00ef0611";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"fffd0611";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"11000608";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"060c9204";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"00b80611";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"ffee0611";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"0b00e804";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"003f0611";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"ff4e0611";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"06f9a104";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"ff690611";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"09003b04";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"00510611";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"ff8f0611";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"03018638";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"03ff4710";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"00facd04";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"00250705";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"11033504";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"ff630705";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"15fa7f04";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"00480705";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"ff810705";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"16040018";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"0c02f910";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"04044d08";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"00fc7f04";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"00150705";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"ff630705";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"18006004";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"005b0705";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"ff6f0705";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"1001eb04";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"ff860705";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"01170705";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"0700e708";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"04043804";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"ff780705";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"00500705";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"11000004";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"ffac0705";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"01990705";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"0205d934";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"0307f820";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"04fae410";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"00fc9808";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"02ff5e04";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"ffa30705";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"00ca0705";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"09004b04";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"ff670705";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"00310705";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"0d008008";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"0f006804";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"00910705";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"fff10705";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"0303b804";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"ffff0705";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"00b40705";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"050e1d0c";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"06105808";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"14004f04";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"00a50705";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"ffd30705";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"ff9c0705";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"0f006f04";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"003a0705";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"ff840705";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"06f84104";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"ff6a0705";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"0c008608";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"0207e904";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"00700705";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"fff50705";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"ff9b0705";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"03018628";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"03fea808";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"00facd04";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"003807dd";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"ff6207dd";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"15f7030c";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"0f007404";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"ff8a07dd";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"02fb9004";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"016007dd";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"003307dd";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"0b00fa0c";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"1af8f804";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"007707dd";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"1e028204";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"ff7507dd";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"ffcb07dd";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"04041d04";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"ff9407dd";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"011807dd";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"0207e93c";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"0304e120";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"05ff8410";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"0e002b08";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"1e026404";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"ffb407dd";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"00ca07dd";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"12004d04";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"ff9b07dd";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"006e07dd";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"03043708";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"04004804";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"ff6707dd";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"fffe07dd";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"04fb4b04";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"007807dd";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"ff9307dd";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"050e1d10";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"060e9008";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"1e023d04";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"ffb807dd";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"007707dd";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"030ebc04";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"ffa607dd";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"007607dd";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"030c5004";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"ff7d07dd";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"05157904";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"007a07dd";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"ffa807dd";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"06fca304";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"ff6e07dd";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"ffea07dd";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"03008128";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"03fea808";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"00facd04";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"003b08b9";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"ff6308b9";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"1af8f804";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"008708b9";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"10001410";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"04043808";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"16040004";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"002308b9";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"ff7908b9";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"0b00d404";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"ff9d08b9";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"00f508b9";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"01fba504";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"002108b9";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"02fa1204";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"ffde08b9";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"ff6608b9";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"01ffcd2c";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"0307f814";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"060e9010";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"08004508";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"16040004";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"ffe508b9";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"00b608b9";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"1703fd04";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"006308b9";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"ffcf08b9";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"ff7808b9";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"060a4e08";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"1e023d04";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"ffd008b9";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"00b708b9";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"02ffe408";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"0f007504";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"001008b9";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"00a308b9";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"0c006404";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"ffce08b9";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"ff3708b9";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"030c5010";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"0800550c";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"1e028708";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"15f6f504";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"ffee08b9";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"ff6108b9";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"000308b9";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"000708b9";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"04e87804";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"ff8108b9";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"00000904";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"00b108b9";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"fff208b9";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"03008124";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"03fea808";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"00facd04";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"003a095d";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"ff64095d";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"1af8f804";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"0074095d";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"0a001910";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"04043808";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"15f70304";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"002f095d";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"ff76095d";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"0b00df04";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"ff8d095d";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"00f1095d";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"1f028704";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"ff68095d";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"002e095d";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"0207e928";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"03036810";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"0500770c";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"0a000404";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"ff6a095d";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"0a000b04";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"00fd095d";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"000b095d";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"ff70095d";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"050e1d10";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"0307f808";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"1d028404";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"003b095d";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"ff97095d";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"060a4e04";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"00a1095d";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"0034095d";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"030c5004";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"ff85095d";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"0013095d";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"06fca304";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"ff75095d";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"ffec095d";
		wait for Clk_period;
		Addr <=  "0001001010111";
		Trees_din <= x"03008128";
		wait for Clk_period;
		Addr <=  "0001001011000";
		Trees_din <= x"03fea808";
		wait for Clk_period;
		Addr <=  "0001001011001";
		Trees_din <= x"00facd04";
		wait for Clk_period;
		Addr <=  "0001001011010";
		Trees_din <= x"003d0a31";
		wait for Clk_period;
		Addr <=  "0001001011011";
		Trees_din <= x"ff650a31";
		wait for Clk_period;
		Addr <=  "0001001011100";
		Trees_din <= x"0b00df08";
		wait for Clk_period;
		Addr <=  "0001001011101";
		Trees_din <= x"03fec304";
		wait for Clk_period;
		Addr <=  "0001001011110";
		Trees_din <= x"00880a31";
		wait for Clk_period;
		Addr <=  "0001001011111";
		Trees_din <= x"ff6a0a31";
		wait for Clk_period;
		Addr <=  "0001001100000";
		Trees_din <= x"04043808";
		wait for Clk_period;
		Addr <=  "0001001100001";
		Trees_din <= x"10021204";
		wait for Clk_period;
		Addr <=  "0001001100010";
		Trees_din <= x"ff760a31";
		wait for Clk_period;
		Addr <=  "0001001100011";
		Trees_din <= x"003b0a31";
		wait for Clk_period;
		Addr <=  "0001001100100";
		Trees_din <= x"0a001408";
		wait for Clk_period;
		Addr <=  "0001001100101";
		Trees_din <= x"08004004";
		wait for Clk_period;
		Addr <=  "0001001100110";
		Trees_din <= x"00040a31";
		wait for Clk_period;
		Addr <=  "0001001100111";
		Trees_din <= x"010b0a31";
		wait for Clk_period;
		Addr <=  "0001001101000";
		Trees_din <= x"1c028504";
		wait for Clk_period;
		Addr <=  "0001001101001";
		Trees_din <= x"ff930a31";
		wait for Clk_period;
		Addr <=  "0001001101010";
		Trees_din <= x"00320a31";
		wait for Clk_period;
		Addr <=  "0001001101011";
		Trees_din <= x"01ffcd24";
		wait for Clk_period;
		Addr <=  "0001001101100";
		Trees_din <= x"0d00b720";
		wait for Clk_period;
		Addr <=  "0001001101101";
		Trees_din <= x"0f007510";
		wait for Clk_period;
		Addr <=  "0001001101110";
		Trees_din <= x"03028a08";
		wait for Clk_period;
		Addr <=  "0001001101111";
		Trees_din <= x"11016e04";
		wait for Clk_period;
		Addr <=  "0001001110000";
		Trees_din <= x"ff700a31";
		wait for Clk_period;
		Addr <=  "0001001110001";
		Trees_din <= x"003d0a31";
		wait for Clk_period;
		Addr <=  "0001001110010";
		Trees_din <= x"0f006b04";
		wait for Clk_period;
		Addr <=  "0001001110011";
		Trees_din <= x"00680a31";
		wait for Clk_period;
		Addr <=  "0001001110100";
		Trees_din <= x"ffe40a31";
		wait for Clk_period;
		Addr <=  "0001001110101";
		Trees_din <= x"1d028608";
		wait for Clk_period;
		Addr <=  "0001001110110";
		Trees_din <= x"060d4204";
		wait for Clk_period;
		Addr <=  "0001001110111";
		Trees_din <= x"005f0a31";
		wait for Clk_period;
		Addr <=  "0001001111000";
		Trees_din <= x"ffe40a31";
		wait for Clk_period;
		Addr <=  "0001001111001";
		Trees_din <= x"0307f804";
		wait for Clk_period;
		Addr <=  "0001001111010";
		Trees_din <= x"ff740a31";
		wait for Clk_period;
		Addr <=  "0001001111011";
		Trees_din <= x"00310a31";
		wait for Clk_period;
		Addr <=  "0001001111100";
		Trees_din <= x"ff580a31";
		wait for Clk_period;
		Addr <=  "0001001111101";
		Trees_din <= x"030c5014";
		wait for Clk_period;
		Addr <=  "0001001111110";
		Trees_din <= x"1f02820c";
		wait for Clk_period;
		Addr <=  "0001001111111";
		Trees_din <= x"15f70d08";
		wait for Clk_period;
		Addr <=  "0001010000000";
		Trees_din <= x"0e002c04";
		wait for Clk_period;
		Addr <=  "0001010000001";
		Trees_din <= x"00300a31";
		wait for Clk_period;
		Addr <=  "0001010000010";
		Trees_din <= x"ffab0a31";
		wait for Clk_period;
		Addr <=  "0001010000011";
		Trees_din <= x"ff640a31";
		wait for Clk_period;
		Addr <=  "0001010000100";
		Trees_din <= x"04018304";
		wait for Clk_period;
		Addr <=  "0001010000101";
		Trees_din <= x"ffa40a31";
		wait for Clk_period;
		Addr <=  "0001010000110";
		Trees_din <= x"004c0a31";
		wait for Clk_period;
		Addr <=  "0001010000111";
		Trees_din <= x"04e87804";
		wait for Clk_period;
		Addr <=  "0001010001000";
		Trees_din <= x"ff8e0a31";
		wait for Clk_period;
		Addr <=  "0001010001001";
		Trees_din <= x"00000904";
		wait for Clk_period;
		Addr <=  "0001010001010";
		Trees_din <= x"00990a31";
		wait for Clk_period;
		Addr <=  "0001010001011";
		Trees_din <= x"fff40a31";
		wait for Clk_period;
		Addr <=  "0001010001100";
		Trees_din <= x"03008120";
		wait for Clk_period;
		Addr <=  "0001010001101";
		Trees_din <= x"03fea808";
		wait for Clk_period;
		Addr <=  "0001010001110";
		Trees_din <= x"00facd04";
		wait for Clk_period;
		Addr <=  "0001010001111";
		Trees_din <= x"003c0b0d";
		wait for Clk_period;
		Addr <=  "0001010010000";
		Trees_din <= x"ff660b0d";
		wait for Clk_period;
		Addr <=  "0001010010001";
		Trees_din <= x"1af8f804";
		wait for Clk_period;
		Addr <=  "0001010010010";
		Trees_din <= x"00750b0d";
		wait for Clk_period;
		Addr <=  "0001010010011";
		Trees_din <= x"0a00190c";
		wait for Clk_period;
		Addr <=  "0001010010100";
		Trees_din <= x"02fa8004";
		wait for Clk_period;
		Addr <=  "0001010010101";
		Trees_din <= x"00c20b0d";
		wait for Clk_period;
		Addr <=  "0001010010110";
		Trees_din <= x"04043804";
		wait for Clk_period;
		Addr <=  "0001010010111";
		Trees_din <= x"ff7b0b0d";
		wait for Clk_period;
		Addr <=  "0001010011000";
		Trees_din <= x"00260b0d";
		wait for Clk_period;
		Addr <=  "0001010011001";
		Trees_din <= x"1f028704";
		wait for Clk_period;
		Addr <=  "0001010011010";
		Trees_din <= x"ff6c0b0d";
		wait for Clk_period;
		Addr <=  "0001010011011";
		Trees_din <= x"002e0b0d";
		wait for Clk_period;
		Addr <=  "0001010011100";
		Trees_din <= x"0001e040";
		wait for Clk_period;
		Addr <=  "0001010011101";
		Trees_din <= x"03067c20";
		wait for Clk_period;
		Addr <=  "0001010011110";
		Trees_din <= x"0500a710";
		wait for Clk_period;
		Addr <=  "0001010011111";
		Trees_din <= x"09004708";
		wait for Clk_period;
		Addr <=  "0001010100000";
		Trees_din <= x"08004004";
		wait for Clk_period;
		Addr <=  "0001010100001";
		Trees_din <= x"ffdb0b0d";
		wait for Clk_period;
		Addr <=  "0001010100010";
		Trees_din <= x"00520b0d";
		wait for Clk_period;
		Addr <=  "0001010100011";
		Trees_din <= x"0a01c304";
		wait for Clk_period;
		Addr <=  "0001010100100";
		Trees_din <= x"ff4f0b0d";
		wait for Clk_period;
		Addr <=  "0001010100101";
		Trees_din <= x"00270b0d";
		wait for Clk_period;
		Addr <=  "0001010100110";
		Trees_din <= x"03043708";
		wait for Clk_period;
		Addr <=  "0001010100111";
		Trees_din <= x"09004904";
		wait for Clk_period;
		Addr <=  "0001010101000";
		Trees_din <= x"ff6c0b0d";
		wait for Clk_period;
		Addr <=  "0001010101001";
		Trees_din <= x"00170b0d";
		wait for Clk_period;
		Addr <=  "0001010101010";
		Trees_din <= x"05043c04";
		wait for Clk_period;
		Addr <=  "0001010101011";
		Trees_din <= x"00460b0d";
		wait for Clk_period;
		Addr <=  "0001010101100";
		Trees_din <= x"ff860b0d";
		wait for Clk_period;
		Addr <=  "0001010101101";
		Trees_din <= x"02fef010";
		wait for Clk_period;
		Addr <=  "0001010101110";
		Trees_din <= x"0c00a208";
		wait for Clk_period;
		Addr <=  "0001010101111";
		Trees_din <= x"1c025104";
		wait for Clk_period;
		Addr <=  "0001010110000";
		Trees_din <= x"006f0b0d";
		wait for Clk_period;
		Addr <=  "0001010110001";
		Trees_din <= x"ffcc0b0d";
		wait for Clk_period;
		Addr <=  "0001010110010";
		Trees_din <= x"10023d04";
		wait for Clk_period;
		Addr <=  "0001010110011";
		Trees_din <= x"00a90b0d";
		wait for Clk_period;
		Addr <=  "0001010110100";
		Trees_din <= x"00070b0d";
		wait for Clk_period;
		Addr <=  "0001010110101";
		Trees_din <= x"0b00e808";
		wait for Clk_period;
		Addr <=  "0001010110110";
		Trees_din <= x"09004704";
		wait for Clk_period;
		Addr <=  "0001010110111";
		Trees_din <= x"004d0b0d";
		wait for Clk_period;
		Addr <=  "0001010111000";
		Trees_din <= x"ff970b0d";
		wait for Clk_period;
		Addr <=  "0001010111001";
		Trees_din <= x"04f84d04";
		wait for Clk_period;
		Addr <=  "0001010111010";
		Trees_din <= x"00340b0d";
		wait for Clk_period;
		Addr <=  "0001010111011";
		Trees_din <= x"ff3e0b0d";
		wait for Clk_period;
		Addr <=  "0001010111100";
		Trees_din <= x"1703fe08";
		wait for Clk_period;
		Addr <=  "0001010111101";
		Trees_din <= x"0e002304";
		wait for Clk_period;
		Addr <=  "0001010111110";
		Trees_din <= x"ffe30b0d";
		wait for Clk_period;
		Addr <=  "0001010111111";
		Trees_din <= x"ff6b0b0d";
		wait for Clk_period;
		Addr <=  "0001011000000";
		Trees_din <= x"0c000c04";
		wait for Clk_period;
		Addr <=  "0001011000001";
		Trees_din <= x"ffa70b0d";
		wait for Clk_period;
		Addr <=  "0001011000010";
		Trees_din <= x"00600b0d";
		wait for Clk_period;
		Addr <=  "0001011000011";
		Trees_din <= x"03ff4714";
		wait for Clk_period;
		Addr <=  "0001011000100";
		Trees_din <= x"00facd04";
		wait for Clk_period;
		Addr <=  "0001011000101";
		Trees_din <= x"00330ba9";
		wait for Clk_period;
		Addr <=  "0001011000110";
		Trees_din <= x"1103350c";
		wait for Clk_period;
		Addr <=  "0001011000111";
		Trees_din <= x"15f70308";
		wait for Clk_period;
		Addr <=  "0001011001000";
		Trees_din <= x"11000204";
		wait for Clk_period;
		Addr <=  "0001011001001";
		Trees_din <= x"ff860ba9";
		wait for Clk_period;
		Addr <=  "0001011001010";
		Trees_din <= x"002d0ba9";
		wait for Clk_period;
		Addr <=  "0001011001011";
		Trees_din <= x"ff660ba9";
		wait for Clk_period;
		Addr <=  "0001011001100";
		Trees_din <= x"00040ba9";
		wait for Clk_period;
		Addr <=  "0001011001101";
		Trees_din <= x"03028a20";
		wait for Clk_period;
		Addr <=  "0001011001110";
		Trees_din <= x"12004510";
		wait for Clk_period;
		Addr <=  "0001011001111";
		Trees_din <= x"05ff4d0c";
		wait for Clk_period;
		Addr <=  "0001011010000";
		Trees_din <= x"14003004";
		wait for Clk_period;
		Addr <=  "0001011010001";
		Trees_din <= x"ff7f0ba9";
		wait for Clk_period;
		Addr <=  "0001011010010";
		Trees_din <= x"09003304";
		wait for Clk_period;
		Addr <=  "0001011010011";
		Trees_din <= x"01270ba9";
		wait for Clk_period;
		Addr <=  "0001011010100";
		Trees_din <= x"003a0ba9";
		wait for Clk_period;
		Addr <=  "0001011010101";
		Trees_din <= x"ff780ba9";
		wait for Clk_period;
		Addr <=  "0001011010110";
		Trees_din <= x"00fcc208";
		wait for Clk_period;
		Addr <=  "0001011010111";
		Trees_din <= x"00fc6b04";
		wait for Clk_period;
		Addr <=  "0001011011000";
		Trees_din <= x"ff9e0ba9";
		wait for Clk_period;
		Addr <=  "0001011011001";
		Trees_din <= x"00d30ba9";
		wait for Clk_period;
		Addr <=  "0001011011010";
		Trees_din <= x"04066204";
		wait for Clk_period;
		Addr <=  "0001011011011";
		Trees_din <= x"ff6a0ba9";
		wait for Clk_period;
		Addr <=  "0001011011100";
		Trees_din <= x"004a0ba9";
		wait for Clk_period;
		Addr <=  "0001011011101";
		Trees_din <= x"01020b14";
		wait for Clk_period;
		Addr <=  "0001011011110";
		Trees_din <= x"0d00b710";
		wait for Clk_period;
		Addr <=  "0001011011111";
		Trees_din <= x"09004708";
		wait for Clk_period;
		Addr <=  "0001011100000";
		Trees_din <= x"0b00e604";
		wait for Clk_period;
		Addr <=  "0001011100001";
		Trees_din <= x"004b0ba9";
		wait for Clk_period;
		Addr <=  "0001011100010";
		Trees_din <= x"fffb0ba9";
		wait for Clk_period;
		Addr <=  "0001011100011";
		Trees_din <= x"05fd5004";
		wait for Clk_period;
		Addr <=  "0001011100100";
		Trees_din <= x"ff390ba9";
		wait for Clk_period;
		Addr <=  "0001011100101";
		Trees_din <= x"00030ba9";
		wait for Clk_period;
		Addr <=  "0001011100110";
		Trees_din <= x"ff640ba9";
		wait for Clk_period;
		Addr <=  "0001011100111";
		Trees_din <= x"06f9a104";
		wait for Clk_period;
		Addr <=  "0001011101000";
		Trees_din <= x"ff850ba9";
		wait for Clk_period;
		Addr <=  "0001011101001";
		Trees_din <= x"ffdf0ba9";
		wait for Clk_period;
		Addr <=  "0001011101010";
		Trees_din <= x"03ff4714";
		wait for Clk_period;
		Addr <=  "0001011101011";
		Trees_din <= x"00facd04";
		wait for Clk_period;
		Addr <=  "0001011101100";
		Trees_din <= x"00300c65";
		wait for Clk_period;
		Addr <=  "0001011101101";
		Trees_din <= x"1103350c";
		wait for Clk_period;
		Addr <=  "0001011101110";
		Trees_din <= x"15f70308";
		wait for Clk_period;
		Addr <=  "0001011101111";
		Trees_din <= x"04041504";
		wait for Clk_period;
		Addr <=  "0001011110000";
		Trees_din <= x"002d0c65";
		wait for Clk_period;
		Addr <=  "0001011110001";
		Trees_din <= x"ff8a0c65";
		wait for Clk_period;
		Addr <=  "0001011110010";
		Trees_din <= x"ff670c65";
		wait for Clk_period;
		Addr <=  "0001011110011";
		Trees_din <= x"00070c65";
		wait for Clk_period;
		Addr <=  "0001011110100";
		Trees_din <= x"0303d430";
		wait for Clk_period;
		Addr <=  "0001011110101";
		Trees_din <= x"05ff9720";
		wait for Clk_period;
		Addr <=  "0001011110110";
		Trees_din <= x"15f77210";
		wait for Clk_period;
		Addr <=  "0001011110111";
		Trees_din <= x"03ff6308";
		wait for Clk_period;
		Addr <=  "0001011111000";
		Trees_din <= x"04053b04";
		wait for Clk_period;
		Addr <=  "0001011111001";
		Trees_din <= x"00080c65";
		wait for Clk_period;
		Addr <=  "0001011111010";
		Trees_din <= x"00890c65";
		wait for Clk_period;
		Addr <=  "0001011111011";
		Trees_din <= x"0b009a04";
		wait for Clk_period;
		Addr <=  "0001011111100";
		Trees_din <= x"00160c65";
		wait for Clk_period;
		Addr <=  "0001011111101";
		Trees_din <= x"ff650c65";
		wait for Clk_period;
		Addr <=  "0001011111110";
		Trees_din <= x"06084608";
		wait for Clk_period;
		Addr <=  "0001011111111";
		Trees_din <= x"12004004";
		wait for Clk_period;
		Addr <=  "0001100000000";
		Trees_din <= x"ff710c65";
		wait for Clk_period;
		Addr <=  "0001100000001";
		Trees_din <= x"00200c65";
		wait for Clk_period;
		Addr <=  "0001100000010";
		Trees_din <= x"0b00b004";
		wait for Clk_period;
		Addr <=  "0001100000011";
		Trees_din <= x"ffdc0c65";
		wait for Clk_period;
		Addr <=  "0001100000100";
		Trees_din <= x"00910c65";
		wait for Clk_period;
		Addr <=  "0001100000101";
		Trees_din <= x"15f76c0c";
		wait for Clk_period;
		Addr <=  "0001100000110";
		Trees_din <= x"09003e04";
		wait for Clk_period;
		Addr <=  "0001100000111";
		Trees_din <= x"ff8b0c65";
		wait for Clk_period;
		Addr <=  "0001100001000";
		Trees_din <= x"00fd9804";
		wait for Clk_period;
		Addr <=  "0001100001001";
		Trees_din <= x"00b90c65";
		wait for Clk_period;
		Addr <=  "0001100001010";
		Trees_din <= x"ffaf0c65";
		wait for Clk_period;
		Addr <=  "0001100001011";
		Trees_din <= x"ff6d0c65";
		wait for Clk_period;
		Addr <=  "0001100001100";
		Trees_din <= x"01020b14";
		wait for Clk_period;
		Addr <=  "0001100001101";
		Trees_din <= x"05fbb604";
		wait for Clk_period;
		Addr <=  "0001100001110";
		Trees_din <= x"ff5e0c65";
		wait for Clk_period;
		Addr <=  "0001100001111";
		Trees_din <= x"0d008108";
		wait for Clk_period;
		Addr <=  "0001100010000";
		Trees_din <= x"14003c04";
		wait for Clk_period;
		Addr <=  "0001100010001";
		Trees_din <= x"ffcf0c65";
		wait for Clk_period;
		Addr <=  "0001100010010";
		Trees_din <= x"00370c65";
		wait for Clk_period;
		Addr <=  "0001100010011";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "0001100010100";
		Trees_din <= x"ff9e0c65";
		wait for Clk_period;
		Addr <=  "0001100010101";
		Trees_din <= x"00750c65";
		wait for Clk_period;
		Addr <=  "0001100010110";
		Trees_din <= x"06f9a104";
		wait for Clk_period;
		Addr <=  "0001100010111";
		Trees_din <= x"ff8c0c65";
		wait for Clk_period;
		Addr <=  "0001100011000";
		Trees_din <= x"ffe30c65";
		wait for Clk_period;
		Addr <=  "0001100011001";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0001100011010";
		Trees_din <= x"03fea808";
		wait for Clk_period;
		Addr <=  "0001100011011";
		Trees_din <= x"00facd04";
		wait for Clk_period;
		Addr <=  "0001100011100";
		Trees_din <= x"00380d1d";
		wait for Clk_period;
		Addr <=  "0001100011101";
		Trees_din <= x"ff680d1d";
		wait for Clk_period;
		Addr <=  "0001100011110";
		Trees_din <= x"03028a24";
		wait for Clk_period;
		Addr <=  "0001100011111";
		Trees_din <= x"04015d0c";
		wait for Clk_period;
		Addr <=  "0001100100000";
		Trees_din <= x"0c02d804";
		wait for Clk_period;
		Addr <=  "0001100100001";
		Trees_din <= x"ff710d1d";
		wait for Clk_period;
		Addr <=  "0001100100010";
		Trees_din <= x"0e002604";
		wait for Clk_period;
		Addr <=  "0001100100011";
		Trees_din <= x"00ad0d1d";
		wait for Clk_period;
		Addr <=  "0001100100100";
		Trees_din <= x"ffab0d1d";
		wait for Clk_period;
		Addr <=  "0001100100101";
		Trees_din <= x"1b02440c";
		wait for Clk_period;
		Addr <=  "0001100100110";
		Trees_din <= x"1e023d04";
		wait for Clk_period;
		Addr <=  "0001100100111";
		Trees_din <= x"ffa40d1d";
		wait for Clk_period;
		Addr <=  "0001100101000";
		Trees_din <= x"1e060004";
		wait for Clk_period;
		Addr <=  "0001100101001";
		Trees_din <= x"00f90d1d";
		wait for Clk_period;
		Addr <=  "0001100101010";
		Trees_din <= x"fff50d1d";
		wait for Clk_period;
		Addr <=  "0001100101011";
		Trees_din <= x"04018304";
		wait for Clk_period;
		Addr <=  "0001100101100";
		Trees_din <= x"00ba0d1d";
		wait for Clk_period;
		Addr <=  "0001100101101";
		Trees_din <= x"0b00d104";
		wait for Clk_period;
		Addr <=  "0001100101110";
		Trees_din <= x"ff860d1d";
		wait for Clk_period;
		Addr <=  "0001100101111";
		Trees_din <= x"000d0d1d";
		wait for Clk_period;
		Addr <=  "0001100110000";
		Trees_din <= x"0c018720";
		wait for Clk_period;
		Addr <=  "0001100110001";
		Trees_din <= x"1703bf10";
		wait for Clk_period;
		Addr <=  "0001100110010";
		Trees_din <= x"1100d708";
		wait for Clk_period;
		Addr <=  "0001100110011";
		Trees_din <= x"11000804";
		wait for Clk_period;
		Addr <=  "0001100110100";
		Trees_din <= x"ffff0d1d";
		wait for Clk_period;
		Addr <=  "0001100110101";
		Trees_din <= x"ff710d1d";
		wait for Clk_period;
		Addr <=  "0001100110110";
		Trees_din <= x"05fe2d04";
		wait for Clk_period;
		Addr <=  "0001100110111";
		Trees_din <= x"00ab0d1d";
		wait for Clk_period;
		Addr <=  "0001100111000";
		Trees_din <= x"002d0d1d";
		wait for Clk_period;
		Addr <=  "0001100111001";
		Trees_din <= x"0a00b508";
		wait for Clk_period;
		Addr <=  "0001100111010";
		Trees_din <= x"04032504";
		wait for Clk_period;
		Addr <=  "0001100111011";
		Trees_din <= x"00190d1d";
		wait for Clk_period;
		Addr <=  "0001100111100";
		Trees_din <= x"ff850d1d";
		wait for Clk_period;
		Addr <=  "0001100111101";
		Trees_din <= x"09003f04";
		wait for Clk_period;
		Addr <=  "0001100111110";
		Trees_din <= x"00da0d1d";
		wait for Clk_period;
		Addr <=  "0001100111111";
		Trees_din <= x"00230d1d";
		wait for Clk_period;
		Addr <=  "0001101000000";
		Trees_din <= x"00008e0c";
		wait for Clk_period;
		Addr <=  "0001101000001";
		Trees_din <= x"0e004a08";
		wait for Clk_period;
		Addr <=  "0001101000010";
		Trees_din <= x"11017804";
		wait for Clk_period;
		Addr <=  "0001101000011";
		Trees_din <= x"006e0d1d";
		wait for Clk_period;
		Addr <=  "0001101000100";
		Trees_din <= x"ffcf0d1d";
		wait for Clk_period;
		Addr <=  "0001101000101";
		Trees_din <= x"ffa60d1d";
		wait for Clk_period;
		Addr <=  "0001101000110";
		Trees_din <= x"ff9a0d1d";
		wait for Clk_period;
		Addr <=  "0001101000111";
		Trees_din <= x"03fea808";
		wait for Clk_period;
		Addr <=  "0001101001000";
		Trees_din <= x"00facd04";
		wait for Clk_period;
		Addr <=  "0001101001001";
		Trees_din <= x"00360db9";
		wait for Clk_period;
		Addr <=  "0001101001010";
		Trees_din <= x"ff690db9";
		wait for Clk_period;
		Addr <=  "0001101001011";
		Trees_din <= x"0307f818";
		wait for Clk_period;
		Addr <=  "0001101001100";
		Trees_din <= x"08005b14";
		wait for Clk_period;
		Addr <=  "0001101001101";
		Trees_din <= x"08005610";
		wait for Clk_period;
		Addr <=  "0001101001110";
		Trees_din <= x"0d007908";
		wait for Clk_period;
		Addr <=  "0001101001111";
		Trees_din <= x"0e003304";
		wait for Clk_period;
		Addr <=  "0001101010000";
		Trees_din <= x"ffb50db9";
		wait for Clk_period;
		Addr <=  "0001101010001";
		Trees_din <= x"000b0db9";
		wait for Clk_period;
		Addr <=  "0001101010010";
		Trees_din <= x"00fd9404";
		wait for Clk_period;
		Addr <=  "0001101010011";
		Trees_din <= x"00640db9";
		wait for Clk_period;
		Addr <=  "0001101010100";
		Trees_din <= x"fff20db9";
		wait for Clk_period;
		Addr <=  "0001101010101";
		Trees_din <= x"ff6d0db9";
		wait for Clk_period;
		Addr <=  "0001101010110";
		Trees_din <= x"009f0db9";
		wait for Clk_period;
		Addr <=  "0001101010111";
		Trees_din <= x"0200051c";
		wait for Clk_period;
		Addr <=  "0001101011000";
		Trees_din <= x"0f007510";
		wait for Clk_period;
		Addr <=  "0001101011001";
		Trees_din <= x"0f007008";
		wait for Clk_period;
		Addr <=  "0001101011010";
		Trees_din <= x"0e004904";
		wait for Clk_period;
		Addr <=  "0001101011011";
		Trees_din <= x"007a0db9";
		wait for Clk_period;
		Addr <=  "0001101011100";
		Trees_din <= x"ffcc0db9";
		wait for Clk_period;
		Addr <=  "0001101011101";
		Trees_din <= x"0d006d04";
		wait for Clk_period;
		Addr <=  "0001101011110";
		Trees_din <= x"002a0db9";
		wait for Clk_period;
		Addr <=  "0001101011111";
		Trees_din <= x"ff6c0db9";
		wait for Clk_period;
		Addr <=  "0001101100000";
		Trees_din <= x"0a001808";
		wait for Clk_period;
		Addr <=  "0001101100001";
		Trees_din <= x"08004204";
		wait for Clk_period;
		Addr <=  "0001101100010";
		Trees_din <= x"ffe40db9";
		wait for Clk_period;
		Addr <=  "0001101100011";
		Trees_din <= x"00630db9";
		wait for Clk_period;
		Addr <=  "0001101100100";
		Trees_din <= x"00a30db9";
		wait for Clk_period;
		Addr <=  "0001101100101";
		Trees_din <= x"07f9be0c";
		wait for Clk_period;
		Addr <=  "0001101100110";
		Trees_din <= x"0a003408";
		wait for Clk_period;
		Addr <=  "0001101100111";
		Trees_din <= x"050c8504";
		wait for Clk_period;
		Addr <=  "0001101101000";
		Trees_din <= x"00350db9";
		wait for Clk_period;
		Addr <=  "0001101101001";
		Trees_din <= x"ffa50db9";
		wait for Clk_period;
		Addr <=  "0001101101010";
		Trees_din <= x"ff6f0db9";
		wait for Clk_period;
		Addr <=  "0001101101011";
		Trees_din <= x"0f008204";
		wait for Clk_period;
		Addr <=  "0001101101100";
		Trees_din <= x"00710db9";
		wait for Clk_period;
		Addr <=  "0001101101101";
		Trees_din <= x"ffb30db9";
		wait for Clk_period;
		Addr <=  "0001101101110";
		Trees_din <= x"03fea808";
		wait for Clk_period;
		Addr <=  "0001101101111";
		Trees_din <= x"00facd04";
		wait for Clk_period;
		Addr <=  "0001101110000";
		Trees_din <= x"00340e45";
		wait for Clk_period;
		Addr <=  "0001101110001";
		Trees_din <= x"ff690e45";
		wait for Clk_period;
		Addr <=  "0001101110010";
		Trees_din <= x"01ffde28";
		wait for Clk_period;
		Addr <=  "0001101110011";
		Trees_din <= x"0d00ae20";
		wait for Clk_period;
		Addr <=  "0001101110100";
		Trees_din <= x"0f007510";
		wait for Clk_period;
		Addr <=  "0001101110101";
		Trees_din <= x"08003c08";
		wait for Clk_period;
		Addr <=  "0001101110110";
		Trees_din <= x"01fdca04";
		wait for Clk_period;
		Addr <=  "0001101110111";
		Trees_din <= x"ffbf0e45";
		wait for Clk_period;
		Addr <=  "0001101111000";
		Trees_din <= x"00c70e45";
		wait for Clk_period;
		Addr <=  "0001101111001";
		Trees_din <= x"18006b04";
		wait for Clk_period;
		Addr <=  "0001101111010";
		Trees_din <= x"ff5f0e45";
		wait for Clk_period;
		Addr <=  "0001101111011";
		Trees_din <= x"fffd0e45";
		wait for Clk_period;
		Addr <=  "0001101111100";
		Trees_din <= x"0f007808";
		wait for Clk_period;
		Addr <=  "0001101111101";
		Trees_din <= x"11000904";
		wait for Clk_period;
		Addr <=  "0001101111110";
		Trees_din <= x"00e20e45";
		wait for Clk_period;
		Addr <=  "0001101111111";
		Trees_din <= x"001c0e45";
		wait for Clk_period;
		Addr <=  "0001110000000";
		Trees_din <= x"0303b804";
		wait for Clk_period;
		Addr <=  "0001110000001";
		Trees_din <= x"ffe10e45";
		wait for Clk_period;
		Addr <=  "0001110000010";
		Trees_din <= x"00340e45";
		wait for Clk_period;
		Addr <=  "0001110000011";
		Trees_din <= x"04ffd804";
		wait for Clk_period;
		Addr <=  "0001110000100";
		Trees_din <= x"00040e45";
		wait for Clk_period;
		Addr <=  "0001110000101";
		Trees_din <= x"ff6b0e45";
		wait for Clk_period;
		Addr <=  "0001110000110";
		Trees_din <= x"030c5010";
		wait for Clk_period;
		Addr <=  "0001110000111";
		Trees_din <= x"1f028208";
		wait for Clk_period;
		Addr <=  "0001110001000";
		Trees_din <= x"15f6f504";
		wait for Clk_period;
		Addr <=  "0001110001001";
		Trees_din <= x"ffe60e45";
		wait for Clk_period;
		Addr <=  "0001110001010";
		Trees_din <= x"ff710e45";
		wait for Clk_period;
		Addr <=  "0001110001011";
		Trees_din <= x"19000204";
		wait for Clk_period;
		Addr <=  "0001110001100";
		Trees_din <= x"fffe0e45";
		wait for Clk_period;
		Addr <=  "0001110001101";
		Trees_din <= x"fff20e45";
		wait for Clk_period;
		Addr <=  "0001110001110";
		Trees_din <= x"01020b04";
		wait for Clk_period;
		Addr <=  "0001110001111";
		Trees_din <= x"00770e45";
		wait for Clk_period;
		Addr <=  "0001110010000";
		Trees_din <= x"ffd30e45";
		wait for Clk_period;
		Addr <=  "0001110010001";
		Trees_din <= x"03fea808";
		wait for Clk_period;
		Addr <=  "0001110010010";
		Trees_din <= x"00facd04";
		wait for Clk_period;
		Addr <=  "0001110010011";
		Trees_din <= x"00330ec1";
		wait for Clk_period;
		Addr <=  "0001110010100";
		Trees_din <= x"ff6a0ec1";
		wait for Clk_period;
		Addr <=  "0001110010101";
		Trees_din <= x"17040024";
		wait for Clk_period;
		Addr <=  "0001110010110";
		Trees_din <= x"14002504";
		wait for Clk_period;
		Addr <=  "0001110010111";
		Trees_din <= x"ff7e0ec1";
		wait for Clk_period;
		Addr <=  "0001110011000";
		Trees_din <= x"18004810";
		wait for Clk_period;
		Addr <=  "0001110011001";
		Trees_din <= x"09003908";
		wait for Clk_period;
		Addr <=  "0001110011010";
		Trees_din <= x"03040104";
		wait for Clk_period;
		Addr <=  "0001110011011";
		Trees_din <= x"ffb00ec1";
		wait for Clk_period;
		Addr <=  "0001110011100";
		Trees_din <= x"00130ec1";
		wait for Clk_period;
		Addr <=  "0001110011101";
		Trees_din <= x"0d008904";
		wait for Clk_period;
		Addr <=  "0001110011110";
		Trees_din <= x"00e00ec1";
		wait for Clk_period;
		Addr <=  "0001110011111";
		Trees_din <= x"00440ec1";
		wait for Clk_period;
		Addr <=  "0001110100000";
		Trees_din <= x"0a018208";
		wait for Clk_period;
		Addr <=  "0001110100001";
		Trees_din <= x"1300c504";
		wait for Clk_period;
		Addr <=  "0001110100010";
		Trees_din <= x"00220ec1";
		wait for Clk_period;
		Addr <=  "0001110100011";
		Trees_din <= x"ffc00ec1";
		wait for Clk_period;
		Addr <=  "0001110100100";
		Trees_din <= x"1e028704";
		wait for Clk_period;
		Addr <=  "0001110100101";
		Trees_din <= x"ffab0ec1";
		wait for Clk_period;
		Addr <=  "0001110100110";
		Trees_din <= x"00890ec1";
		wait for Clk_period;
		Addr <=  "0001110100111";
		Trees_din <= x"02fc7304";
		wait for Clk_period;
		Addr <=  "0001110101000";
		Trees_din <= x"ff640ec1";
		wait for Clk_period;
		Addr <=  "0001110101001";
		Trees_din <= x"1e024704";
		wait for Clk_period;
		Addr <=  "0001110101010";
		Trees_din <= x"ff900ec1";
		wait for Clk_period;
		Addr <=  "0001110101011";
		Trees_din <= x"00fe9108";
		wait for Clk_period;
		Addr <=  "0001110101100";
		Trees_din <= x"12004f04";
		wait for Clk_period;
		Addr <=  "0001110101101";
		Trees_din <= x"00140ec1";
		wait for Clk_period;
		Addr <=  "0001110101110";
		Trees_din <= x"00910ec1";
		wait for Clk_period;
		Addr <=  "0001110101111";
		Trees_din <= x"ffc40ec1";
		wait for Clk_period;
		Addr <=  "0001110110000";
		Trees_din <= x"03fea808";
		wait for Clk_period;
		Addr <=  "0001110110001";
		Trees_din <= x"00facd04";
		wait for Clk_period;
		Addr <=  "0001110110010";
		Trees_din <= x"00310f3d";
		wait for Clk_period;
		Addr <=  "0001110110011";
		Trees_din <= x"ff6b0f3d";
		wait for Clk_period;
		Addr <=  "0001110110100";
		Trees_din <= x"01ffde24";
		wait for Clk_period;
		Addr <=  "0001110110101";
		Trees_din <= x"0d00b720";
		wait for Clk_period;
		Addr <=  "0001110110110";
		Trees_din <= x"0d007910";
		wait for Clk_period;
		Addr <=  "0001110110111";
		Trees_din <= x"10027008";
		wait for Clk_period;
		Addr <=  "0001110111000";
		Trees_din <= x"16033804";
		wait for Clk_period;
		Addr <=  "0001110111001";
		Trees_din <= x"00820f3d";
		wait for Clk_period;
		Addr <=  "0001110111010";
		Trees_din <= x"fff60f3d";
		wait for Clk_period;
		Addr <=  "0001110111011";
		Trees_din <= x"03079404";
		wait for Clk_period;
		Addr <=  "0001110111100";
		Trees_din <= x"ff650f3d";
		wait for Clk_period;
		Addr <=  "0001110111101";
		Trees_din <= x"00150f3d";
		wait for Clk_period;
		Addr <=  "0001110111110";
		Trees_din <= x"07ff1e08";
		wait for Clk_period;
		Addr <=  "0001110111111";
		Trees_din <= x"0d008604";
		wait for Clk_period;
		Addr <=  "0001111000000";
		Trees_din <= x"00740f3d";
		wait for Clk_period;
		Addr <=  "0001111000001";
		Trees_din <= x"000d0f3d";
		wait for Clk_period;
		Addr <=  "0001111000010";
		Trees_din <= x"1b024804";
		wait for Clk_period;
		Addr <=  "0001111000011";
		Trees_din <= x"005e0f3d";
		wait for Clk_period;
		Addr <=  "0001111000100";
		Trees_din <= x"ffa90f3d";
		wait for Clk_period;
		Addr <=  "0001111000101";
		Trees_din <= x"ff7f0f3d";
		wait for Clk_period;
		Addr <=  "0001111000110";
		Trees_din <= x"030c500c";
		wait for Clk_period;
		Addr <=  "0001111000111";
		Trees_din <= x"1f028208";
		wait for Clk_period;
		Addr <=  "0001111001000";
		Trees_din <= x"16040004";
		wait for Clk_period;
		Addr <=  "0001111001001";
		Trees_din <= x"ff710f3d";
		wait for Clk_period;
		Addr <=  "0001111001010";
		Trees_din <= x"ffd30f3d";
		wait for Clk_period;
		Addr <=  "0001111001011";
		Trees_din <= x"fff50f3d";
		wait for Clk_period;
		Addr <=  "0001111001100";
		Trees_din <= x"01020b04";
		wait for Clk_period;
		Addr <=  "0001111001101";
		Trees_din <= x"006e0f3d";
		wait for Clk_period;
		Addr <=  "0001111001110";
		Trees_din <= x"ffda0f3d";
		wait for Clk_period;
		Addr <=  "0001111001111";
		Trees_din <= x"03fea808";
		wait for Clk_period;
		Addr <=  "0001111010000";
		Trees_din <= x"00facd04";
		wait for Clk_period;
		Addr <=  "0001111010001";
		Trees_din <= x"00300fe1";
		wait for Clk_period;
		Addr <=  "0001111010010";
		Trees_din <= x"ff6c0fe1";
		wait for Clk_period;
		Addr <=  "0001111010011";
		Trees_din <= x"1e025f2c";
		wait for Clk_period;
		Addr <=  "0001111010100";
		Trees_din <= x"12004d10";
		wait for Clk_period;
		Addr <=  "0001111010101";
		Trees_din <= x"030cf40c";
		wait for Clk_period;
		Addr <=  "0001111010110";
		Trees_din <= x"06f9a104";
		wait for Clk_period;
		Addr <=  "0001111010111";
		Trees_din <= x"00610fe1";
		wait for Clk_period;
		Addr <=  "0001111011000";
		Trees_din <= x"1d025404";
		wait for Clk_period;
		Addr <=  "0001111011001";
		Trees_din <= x"ffd70fe1";
		wait for Clk_period;
		Addr <=  "0001111011010";
		Trees_din <= x"ff500fe1";
		wait for Clk_period;
		Addr <=  "0001111011011";
		Trees_din <= x"00580fe1";
		wait for Clk_period;
		Addr <=  "0001111011100";
		Trees_din <= x"11000210";
		wait for Clk_period;
		Addr <=  "0001111011101";
		Trees_din <= x"0b00df08";
		wait for Clk_period;
		Addr <=  "0001111011110";
		Trees_din <= x"1e025204";
		wait for Clk_period;
		Addr <=  "0001111011111";
		Trees_din <= x"ff730fe1";
		wait for Clk_period;
		Addr <=  "0001111100000";
		Trees_din <= x"00050fe1";
		wait for Clk_period;
		Addr <=  "0001111100001";
		Trees_din <= x"07002504";
		wait for Clk_period;
		Addr <=  "0001111100010";
		Trees_din <= x"00000fe1";
		wait for Clk_period;
		Addr <=  "0001111100011";
		Trees_din <= x"00750fe1";
		wait for Clk_period;
		Addr <=  "0001111100100";
		Trees_din <= x"18008808";
		wait for Clk_period;
		Addr <=  "0001111100101";
		Trees_din <= x"16040004";
		wait for Clk_period;
		Addr <=  "0001111100110";
		Trees_din <= x"004f0fe1";
		wait for Clk_period;
		Addr <=  "0001111100111";
		Trees_din <= x"00f80fe1";
		wait for Clk_period;
		Addr <=  "0001111101000";
		Trees_din <= x"ffc70fe1";
		wait for Clk_period;
		Addr <=  "0001111101001";
		Trees_din <= x"10000908";
		wait for Clk_period;
		Addr <=  "0001111101010";
		Trees_din <= x"00fe5d04";
		wait for Clk_period;
		Addr <=  "0001111101011";
		Trees_din <= x"00c40fe1";
		wait for Clk_period;
		Addr <=  "0001111101100";
		Trees_din <= x"000e0fe1";
		wait for Clk_period;
		Addr <=  "0001111101101";
		Trees_din <= x"1703ff10";
		wait for Clk_period;
		Addr <=  "0001111101110";
		Trees_din <= x"0306ca08";
		wait for Clk_period;
		Addr <=  "0001111101111";
		Trees_din <= x"0500e804";
		wait for Clk_period;
		Addr <=  "0001111110000";
		Trees_din <= x"00130fe1";
		wait for Clk_period;
		Addr <=  "0001111110001";
		Trees_din <= x"ff9f0fe1";
		wait for Clk_period;
		Addr <=  "0001111110010";
		Trees_din <= x"00fcaa04";
		wait for Clk_period;
		Addr <=  "0001111110011";
		Trees_din <= x"ffc50fe1";
		wait for Clk_period;
		Addr <=  "0001111110100";
		Trees_din <= x"006a0fe1";
		wait for Clk_period;
		Addr <=  "0001111110101";
		Trees_din <= x"01fe7504";
		wait for Clk_period;
		Addr <=  "0001111110110";
		Trees_din <= x"ff730fe1";
		wait for Clk_period;
		Addr <=  "0001111110111";
		Trees_din <= x"fffa0fe1";
		wait for Clk_period;
		Addr <=  "0001111111000";
		Trees_din <= x"03fea808";
		wait for Clk_period;
		Addr <=  "0001111111001";
		Trees_din <= x"00facd04";
		wait for Clk_period;
		Addr <=  "0001111111010";
		Trees_din <= x"002e10ad";
		wait for Clk_period;
		Addr <=  "0001111111011";
		Trees_din <= x"ff6d10ad";
		wait for Clk_period;
		Addr <=  "0001111111100";
		Trees_din <= x"02fef034";
		wait for Clk_period;
		Addr <=  "0001111111101";
		Trees_din <= x"02fdc120";
		wait for Clk_period;
		Addr <=  "0001111111110";
		Trees_din <= x"0d008110";
		wait for Clk_period;
		Addr <=  "0001111111111";
		Trees_din <= x"060a0a08";
		wait for Clk_period;
		Addr <=  "0010000000000";
		Trees_din <= x"0608ee04";
		wait for Clk_period;
		Addr <=  "0010000000001";
		Trees_din <= x"ffeb10ad";
		wait for Clk_period;
		Addr <=  "0010000000010";
		Trees_din <= x"007110ad";
		wait for Clk_period;
		Addr <=  "0010000000011";
		Trees_din <= x"16020204";
		wait for Clk_period;
		Addr <=  "0010000000100";
		Trees_din <= x"00a910ad";
		wait for Clk_period;
		Addr <=  "0010000000101";
		Trees_din <= x"ff9a10ad";
		wait for Clk_period;
		Addr <=  "0010000000110";
		Trees_din <= x"00fd9408";
		wait for Clk_period;
		Addr <=  "0010000000111";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "0010000001000";
		Trees_din <= x"ffc210ad";
		wait for Clk_period;
		Addr <=  "0010000001001";
		Trees_din <= x"009c10ad";
		wait for Clk_period;
		Addr <=  "0010000001010";
		Trees_din <= x"04007504";
		wait for Clk_period;
		Addr <=  "0010000001011";
		Trees_din <= x"004110ad";
		wait for Clk_period;
		Addr <=  "0010000001100";
		Trees_din <= x"ffb810ad";
		wait for Clk_period;
		Addr <=  "0010000001101";
		Trees_din <= x"03021004";
		wait for Clk_period;
		Addr <=  "0010000001110";
		Trees_din <= x"ff9a10ad";
		wait for Clk_period;
		Addr <=  "0010000001111";
		Trees_din <= x"05001308";
		wait for Clk_period;
		Addr <=  "0010000010000";
		Trees_din <= x"1afc7904";
		wait for Clk_period;
		Addr <=  "0010000010001";
		Trees_din <= x"00d110ad";
		wait for Clk_period;
		Addr <=  "0010000010010";
		Trees_din <= x"fffc10ad";
		wait for Clk_period;
		Addr <=  "0010000010011";
		Trees_din <= x"03067c04";
		wait for Clk_period;
		Addr <=  "0010000010100";
		Trees_din <= x"ffb610ad";
		wait for Clk_period;
		Addr <=  "0010000010101";
		Trees_din <= x"005c10ad";
		wait for Clk_period;
		Addr <=  "0010000010110";
		Trees_din <= x"1d025e14";
		wait for Clk_period;
		Addr <=  "0010000010111";
		Trees_din <= x"0201110c";
		wait for Clk_period;
		Addr <=  "0010000011000";
		Trees_din <= x"13009b04";
		wait for Clk_period;
		Addr <=  "0010000011001";
		Trees_din <= x"ffe410ad";
		wait for Clk_period;
		Addr <=  "0010000011010";
		Trees_din <= x"0e003204";
		wait for Clk_period;
		Addr <=  "0010000011011";
		Trees_din <= x"002710ad";
		wait for Clk_period;
		Addr <=  "0010000011100";
		Trees_din <= x"00a710ad";
		wait for Clk_period;
		Addr <=  "0010000011101";
		Trees_din <= x"030c5004";
		wait for Clk_period;
		Addr <=  "0010000011110";
		Trees_din <= x"ff9910ad";
		wait for Clk_period;
		Addr <=  "0010000011111";
		Trees_din <= x"002e10ad";
		wait for Clk_period;
		Addr <=  "0010000100000";
		Trees_din <= x"0d006708";
		wait for Clk_period;
		Addr <=  "0010000100001";
		Trees_din <= x"01fd0104";
		wait for Clk_period;
		Addr <=  "0010000100010";
		Trees_din <= x"006a10ad";
		wait for Clk_period;
		Addr <=  "0010000100011";
		Trees_din <= x"fff610ad";
		wait for Clk_period;
		Addr <=  "0010000100100";
		Trees_din <= x"02015508";
		wait for Clk_period;
		Addr <=  "0010000100101";
		Trees_din <= x"05011c04";
		wait for Clk_period;
		Addr <=  "0010000100110";
		Trees_din <= x"ff4e10ad";
		wait for Clk_period;
		Addr <=  "0010000100111";
		Trees_din <= x"ffeb10ad";
		wait for Clk_period;
		Addr <=  "0010000101000";
		Trees_din <= x"02051804";
		wait for Clk_period;
		Addr <=  "0010000101001";
		Trees_din <= x"002d10ad";
		wait for Clk_period;
		Addr <=  "0010000101010";
		Trees_din <= x"ffa910ad";
		wait for Clk_period;
		Addr <=  "0010000101011";
		Trees_din <= x"03fde504";
		wait for Clk_period;
		Addr <=  "0010000101100";
		Trees_din <= x"ff6f1151";
		wait for Clk_period;
		Addr <=  "0010000101101";
		Trees_din <= x"0900472c";
		wait for Clk_period;
		Addr <=  "0010000101110";
		Trees_din <= x"09004620";
		wait for Clk_period;
		Addr <=  "0010000101111";
		Trees_din <= x"0f007510";
		wait for Clk_period;
		Addr <=  "0010000110000";
		Trees_din <= x"08003c08";
		wait for Clk_period;
		Addr <=  "0010000110001";
		Trees_din <= x"1e026604";
		wait for Clk_period;
		Addr <=  "0010000110010";
		Trees_din <= x"ffa21151";
		wait for Clk_period;
		Addr <=  "0010000110011";
		Trees_din <= x"00881151";
		wait for Clk_period;
		Addr <=  "0010000110100";
		Trees_din <= x"0f006b04";
		wait for Clk_period;
		Addr <=  "0010000110101";
		Trees_din <= x"00121151";
		wait for Clk_period;
		Addr <=  "0010000110110";
		Trees_din <= x"ffa81151";
		wait for Clk_period;
		Addr <=  "0010000110111";
		Trees_din <= x"1603ec08";
		wait for Clk_period;
		Addr <=  "0010000111000";
		Trees_din <= x"1702a604";
		wait for Clk_period;
		Addr <=  "0010000111001";
		Trees_din <= x"003a1151";
		wait for Clk_period;
		Addr <=  "0010000111010";
		Trees_din <= x"ffc51151";
		wait for Clk_period;
		Addr <=  "0010000111011";
		Trees_din <= x"0f007804";
		wait for Clk_period;
		Addr <=  "0010000111100";
		Trees_din <= x"00731151";
		wait for Clk_period;
		Addr <=  "0010000111101";
		Trees_din <= x"00181151";
		wait for Clk_period;
		Addr <=  "0010000111110";
		Trees_din <= x"0b00b108";
		wait for Clk_period;
		Addr <=  "0010000111111";
		Trees_din <= x"1300aa04";
		wait for Clk_period;
		Addr <=  "0010001000000";
		Trees_din <= x"00d61151";
		wait for Clk_period;
		Addr <=  "0010001000001";
		Trees_din <= x"00381151";
		wait for Clk_period;
		Addr <=  "0010001000010";
		Trees_din <= x"ffbf1151";
		wait for Clk_period;
		Addr <=  "0010001000011";
		Trees_din <= x"1900000c";
		wait for Clk_period;
		Addr <=  "0010001000100";
		Trees_din <= x"00fcf104";
		wait for Clk_period;
		Addr <=  "0010001000101";
		Trees_din <= x"ffed1151";
		wait for Clk_period;
		Addr <=  "0010001000110";
		Trees_din <= x"17011f04";
		wait for Clk_period;
		Addr <=  "0010001000111";
		Trees_din <= x"ffef1151";
		wait for Clk_period;
		Addr <=  "0010001001000";
		Trees_din <= x"ff651151";
		wait for Clk_period;
		Addr <=  "0010001001001";
		Trees_din <= x"00fed010";
		wait for Clk_period;
		Addr <=  "0010001001010";
		Trees_din <= x"1e028008";
		wait for Clk_period;
		Addr <=  "0010001001011";
		Trees_din <= x"08004704";
		wait for Clk_period;
		Addr <=  "0010001001100";
		Trees_din <= x"00251151";
		wait for Clk_period;
		Addr <=  "0010001001101";
		Trees_din <= x"ffb11151";
		wait for Clk_period;
		Addr <=  "0010001001110";
		Trees_din <= x"19000204";
		wait for Clk_period;
		Addr <=  "0010001001111";
		Trees_din <= x"00d51151";
		wait for Clk_period;
		Addr <=  "0010001010000";
		Trees_din <= x"00421151";
		wait for Clk_period;
		Addr <=  "0010001010001";
		Trees_din <= x"1b027004";
		wait for Clk_period;
		Addr <=  "0010001010010";
		Trees_din <= x"000b1151";
		wait for Clk_period;
		Addr <=  "0010001010011";
		Trees_din <= x"ff861151";
		wait for Clk_period;
		Addr <=  "0010001010100";
		Trees_din <= x"03fde504";
		wait for Clk_period;
		Addr <=  "0010001010101";
		Trees_din <= x"ff711205";
		wait for Clk_period;
		Addr <=  "0010001010110";
		Trees_din <= x"03008118";
		wait for Clk_period;
		Addr <=  "0010001010111";
		Trees_din <= x"08004714";
		wait for Clk_period;
		Addr <=  "0010001011000";
		Trees_din <= x"08004610";
		wait for Clk_period;
		Addr <=  "0010001011001";
		Trees_din <= x"06068d08";
		wait for Clk_period;
		Addr <=  "0010001011010";
		Trees_din <= x"0e002404";
		wait for Clk_period;
		Addr <=  "0010001011011";
		Trees_din <= x"ffaa1205";
		wait for Clk_period;
		Addr <=  "0010001011100";
		Trees_din <= x"00431205";
		wait for Clk_period;
		Addr <=  "0010001011101";
		Trees_din <= x"0d005f04";
		wait for Clk_period;
		Addr <=  "0010001011110";
		Trees_din <= x"00451205";
		wait for Clk_period;
		Addr <=  "0010001011111";
		Trees_din <= x"ff791205";
		wait for Clk_period;
		Addr <=  "0010001100000";
		Trees_din <= x"00cc1205";
		wait for Clk_period;
		Addr <=  "0010001100001";
		Trees_din <= x"ff7b1205";
		wait for Clk_period;
		Addr <=  "0010001100010";
		Trees_din <= x"09004720";
		wait for Clk_period;
		Addr <=  "0010001100011";
		Trees_din <= x"04036410";
		wait for Clk_period;
		Addr <=  "0010001100100";
		Trees_din <= x"1e026408";
		wait for Clk_period;
		Addr <=  "0010001100101";
		Trees_din <= x"0b00c904";
		wait for Clk_period;
		Addr <=  "0010001100110";
		Trees_din <= x"00311205";
		wait for Clk_period;
		Addr <=  "0010001100111";
		Trees_din <= x"ffc21205";
		wait for Clk_period;
		Addr <=  "0010001101000";
		Trees_din <= x"1000d804";
		wait for Clk_period;
		Addr <=  "0010001101001";
		Trees_din <= x"00591205";
		wait for Clk_period;
		Addr <=  "0010001101010";
		Trees_din <= x"00051205";
		wait for Clk_period;
		Addr <=  "0010001101011";
		Trees_din <= x"09004008";
		wait for Clk_period;
		Addr <=  "0010001101100";
		Trees_din <= x"12003704";
		wait for Clk_period;
		Addr <=  "0010001101101";
		Trees_din <= x"00171205";
		wait for Clk_period;
		Addr <=  "0010001101110";
		Trees_din <= x"ff681205";
		wait for Clk_period;
		Addr <=  "0010001101111";
		Trees_din <= x"1300b304";
		wait for Clk_period;
		Addr <=  "0010001110000";
		Trees_din <= x"ff941205";
		wait for Clk_period;
		Addr <=  "0010001110001";
		Trees_din <= x"00cd1205";
		wait for Clk_period;
		Addr <=  "0010001110010";
		Trees_din <= x"1c028010";
		wait for Clk_period;
		Addr <=  "0010001110011";
		Trees_din <= x"00fd1008";
		wait for Clk_period;
		Addr <=  "0010001110100";
		Trees_din <= x"06093d04";
		wait for Clk_period;
		Addr <=  "0010001110101";
		Trees_din <= x"006e1205";
		wait for Clk_period;
		Addr <=  "0010001110110";
		Trees_din <= x"ffb51205";
		wait for Clk_period;
		Addr <=  "0010001110111";
		Trees_din <= x"03079404";
		wait for Clk_period;
		Addr <=  "0010001111000";
		Trees_din <= x"ff5f1205";
		wait for Clk_period;
		Addr <=  "0010001111001";
		Trees_din <= x"00071205";
		wait for Clk_period;
		Addr <=  "0010001111010";
		Trees_din <= x"02fc7908";
		wait for Clk_period;
		Addr <=  "0010001111011";
		Trees_din <= x"1100a404";
		wait for Clk_period;
		Addr <=  "0010001111100";
		Trees_din <= x"00881205";
		wait for Clk_period;
		Addr <=  "0010001111101";
		Trees_din <= x"fff71205";
		wait for Clk_period;
		Addr <=  "0010001111110";
		Trees_din <= x"0e003d04";
		wait for Clk_period;
		Addr <=  "0010001111111";
		Trees_din <= x"00031205";
		wait for Clk_period;
		Addr <=  "0010010000000";
		Trees_din <= x"ff9d1205";
		wait for Clk_period;
		Addr <=  "0010010000001";
		Trees_din <= x"03fde504";
		wait for Clk_period;
		Addr <=  "0010010000010";
		Trees_din <= x"ff721261";
		wait for Clk_period;
		Addr <=  "0010010000011";
		Trees_din <= x"1701e40c";
		wait for Clk_period;
		Addr <=  "0010010000100";
		Trees_din <= x"1c028808";
		wait for Clk_period;
		Addr <=  "0010010000101";
		Trees_din <= x"03079404";
		wait for Clk_period;
		Addr <=  "0010010000110";
		Trees_din <= x"ff851261";
		wait for Clk_period;
		Addr <=  "0010010000111";
		Trees_din <= x"00391261";
		wait for Clk_period;
		Addr <=  "0010010001000";
		Trees_din <= x"00471261";
		wait for Clk_period;
		Addr <=  "0010010001001";
		Trees_din <= x"17020004";
		wait for Clk_period;
		Addr <=  "0010010001010";
		Trees_din <= x"008b1261";
		wait for Clk_period;
		Addr <=  "0010010001011";
		Trees_din <= x"1b023d0c";
		wait for Clk_period;
		Addr <=  "0010010001100";
		Trees_din <= x"1702f604";
		wait for Clk_period;
		Addr <=  "0010010001101";
		Trees_din <= x"00381261";
		wait for Clk_period;
		Addr <=  "0010010001110";
		Trees_din <= x"01fbe104";
		wait for Clk_period;
		Addr <=  "0010010001111";
		Trees_din <= x"00341261";
		wait for Clk_period;
		Addr <=  "0010010010000";
		Trees_din <= x"ff8e1261";
		wait for Clk_period;
		Addr <=  "0010010010001";
		Trees_din <= x"1d024808";
		wait for Clk_period;
		Addr <=  "0010010010010";
		Trees_din <= x"0d007004";
		wait for Clk_period;
		Addr <=  "0010010010011";
		Trees_din <= x"ffd61261";
		wait for Clk_period;
		Addr <=  "0010010010100";
		Trees_din <= x"007e1261";
		wait for Clk_period;
		Addr <=  "0010010010101";
		Trees_din <= x"0d009a04";
		wait for Clk_period;
		Addr <=  "0010010010110";
		Trees_din <= x"000b1261";
		wait for Clk_period;
		Addr <=  "0010010010111";
		Trees_din <= x"ff8b1261";
		wait for Clk_period;
		Addr <=  "0010010011000";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  3
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"050e1d48";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"0506342c";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"05025514";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"05002d04";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"ff5200a5";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"02fa8408";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"00fdfd04";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"ffa400a5";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"012b00a5";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"0a036704";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"ff5b00a5";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"003700a5";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"02fc160c";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"0700ca08";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"11001d04";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"000000a5";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"026e00a5";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"ff8800a5";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"00fb6004";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"003700a5";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"0b011504";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"ff6e00a5";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"003700a5";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"0202a718";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"13009208";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"01fc5a04";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"003700a5";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"ff8400a5";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"0b00e108";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"19001f04";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"033300a5";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"008900a5";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"00fd2c04";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"ff9000a5";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"017d00a5";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"ff5a00a5";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"02201308";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"07015104";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"047800a5";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"012b00a5";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"ff6f00a5";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"05098550";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"05043c28";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"05025514";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"05002d04";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"ff570179";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"02fa8408";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"12004204";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"01670179";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"ff990179";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"0a036704";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"ff630179";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"00410179";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"02fc0b0c";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"1e027404";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"ff980179";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"07003104";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"01a10179";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"003c0179";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"0d006404";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"00010179";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"ff5e0179";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"07fdba10";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"0b011f0c";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"0b00b408";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"060c1704";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"ff760179";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"00900179";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"ff5f0179";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"00d40179";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"07ffdf08";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"13009804";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"00390179";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"018e0179";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"00fe3d08";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"07013604";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"ff930179";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"01ba0179";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"10001304";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"00290179";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"ff730179";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"02201318";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"07056c14";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"0609450c";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"1e056908";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"09004e04";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"01ad0179";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"006d0179";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"00240179";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"13009204";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"ff7b0179";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"017a0179";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"ffa00179";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"ff670179";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"05063438";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"05025518";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"05002d04";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"ff5b023d";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"02fa8408";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"12004204";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"012e023d";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"ffa1023d";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"03fff508";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"0e004104";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"ff7f023d";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"0070023d";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"ff5d023d";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"02fc160c";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"0700ca08";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"11001d04";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"001b023d";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"0158023d";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"ff92023d";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"01fd780c";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"04ff1c08";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"07ff1704";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"ff70023d";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"001c023d";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"00e3023d";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"0e001a04";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"0023023d";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"ff60023d";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"02201328";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"050e1d10";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"0202a70c";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"0a000304";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"ff83023d";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"0d006304";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"ffc6023d";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"0114023d";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"ff6c023d";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"15f6f908";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"07fb6b04";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"00c8023d";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"ffcb023d";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"08003b08";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"05131704";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"ffe7023d";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"00c5023d";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"1c04ad04";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"013a023d";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"0063023d";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"ff6b023d";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"05063444";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"05025520";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"05002d04";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"ff5e0311";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"02fb1a0c";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"0500c508";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"09003c04";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"00110311";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"013d0311";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"ff8d0311";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"05003908";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"17037804";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"00460311";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"ffad0311";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"01fc3104";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"ffb00311";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"ff600311";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"02fc1610";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"0700ca0c";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"0e003808";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"0f007904";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"ff9f0311";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"00c70311";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"01500311";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"ff990311";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"01fd780c";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"04ff1c08";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"01fb8f04";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"001b0311";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"ff750311";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"00bb0311";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"0e001a04";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"00250311";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"ff650311";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"02201324";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"05157918";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"0203510c";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"030b2708";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"13007804";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"ffe30311";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"00cd0311";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"ff810311";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"06ecd604";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"ff710311";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"03067c04";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"00c70311";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"ffa60311";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"15f6f908";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"0a002904";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"00a30311";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"ffbb0311";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"01020311";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"ff710311";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"0506343c";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"0502551c";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"05002d04";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"ff6003e5";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"02fb1a0c";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"06070104";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"ff9303e5";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"060a7304";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"014903e5";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"ffae03e5";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"05003904";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"ffff03e5";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"01fc3104";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"ffba03e5";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"ff6303e5";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"02fc160c";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"0700ca08";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"14003e04";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"003003e5";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"010a03e5";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"ff9e03e5";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"08004510";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"07fdba08";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"0e001a04";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"003a03e5";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"ff7503e5";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"01fd7804";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"00f103e5";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"ff9503e5";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"ff6a03e5";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"0220132c";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"0513171c";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"02019c0c";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"10033e08";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"08005804";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"00a903e5";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"ff8603e5";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"ff6b03e5";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"0c028008";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"16040004";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"ff5a03e5";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"002503e5";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"0d006d04";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"fff703e5";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"008c03e5";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"15f6f908";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"02051804";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"ff9a03e5";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"00ac03e5";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"07014504";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"00de03e5";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"004903e5";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"ff7803e5";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"05043c2c";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"05002d04";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"ff620489";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"02fbd218";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"01fd330c";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"0401a704";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"ff9f0489";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"00fd0b04";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"001c0489";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"01460489";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"1100a404";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"ff780489";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"1afb4404";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"ffab0489";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"009e0489";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"0503f70c";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"01fc3108";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"03fff504";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"00b50489";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"ff7c0489";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"ff650489";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"00010489";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"05131718";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"0207e914";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"030b2710";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"060d3208";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"07ffa904";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"009b0489";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"00270489";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"09004504";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"ff7e0489";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"005d0489";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"ff770489";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"ff6f0489";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"15f6f908";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"02051804";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"ff9d0489";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"00950489";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"06c00004";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"001d0489";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"00c70489";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"05043c28";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"05002d04";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"ff640525";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"02fbd214";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"01fd330c";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"0401a704";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"ffa50525";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"0606b304";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"00090525";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"01180525";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"1100a404";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"ff7f0525";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"00350525";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"01fceb0c";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"04ff8504";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"ff760525";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"05019e04";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"ff9f0525";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"00ea0525";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"ff680525";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"05157918";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"0207e914";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"030b2710";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"01ff9208";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"00004604";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"00480525";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"ff5c0525";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"09004c04";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"009a0525";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"ffaa0525";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"ff6b0525";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"ff730525";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"15f6f908";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"0d007504";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"007b0525";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"ffab0525";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"06c00004";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"00280525";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"00bc0525";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"0503f724";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"05002d04";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"ff6605b9";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"02fbd214";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"1d027c10";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"09003d08";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"1c027404";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"ff9905b9";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"002505b9";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"0f007804";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"00ec05b9";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"000e05b9";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"ff8f05b9";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"01fc3108";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"03fff504";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"009c05b9";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"ff8705b9";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"ff6a05b9";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"05157918";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"0207e914";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"030b2710";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"1e027008";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"0e002704";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"fff005b9";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"008d05b9";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"0c00c804";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"ff8705b9";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"004005b9";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"ff7305b9";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"ff7805b9";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"15f6f908";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"0d007504";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"006d05b9";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"ffa805b9";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"06c00004";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"002005b9";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"00b105b9";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"05034028";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"05ffaf0c";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"0f005b08";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"00fd7104";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"003e0651";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"ff800651";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"ff650651";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"03fff518";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"01fc3108";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"1703d804";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"00110651";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"01400651";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"0e004108";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"02f9f604";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"00170651";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"ff750651";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"14004b04";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"00cc0651";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"ffeb0651";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"ff6a0651";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"05157918";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"0207e914";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"030b2710";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"07ffdf08";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"01fc0f04";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"ffc00651";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"00650651";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"1300a304";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"ff8d0651";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"003f0651";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"ff7c0651";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"ff7c0651";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"15f71a08";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"07fb6b04";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"00880651";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"ff6f0651";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"00a80651";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"05025524";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"05ffaf0c";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"0f005b08";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"0d005804";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"ff8406dd";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"003d06dd";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"ff6606dd";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"03fff514";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"01fc3108";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"0609a604";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"013106dd";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"000f06dd";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"0e004108";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"02f9f604";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"001906dd";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"ff7a06dd";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"005f06dd";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"ff6f06dd";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"05157918";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"0207e914";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"030b2710";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"09004c08";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"01ffde04";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"001606dd";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"006e06dd";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"0e003c04";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"ff6106dd";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"001406dd";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"ff8606dd";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"ff8006dd";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"15f71a08";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"07fb6b04";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"007c06dd";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"ff7c06dd";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"00a206dd";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"0501c32c";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"05ffaf14";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"0f005b08";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"00fd7104";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"004407a9";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"ff8807a9";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"1f028704";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"ff6507a9";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"1603b904";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"ff7b07a9";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"004207a9";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"03ff8b14";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"0d006e0c";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"13009504";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"ffaf07a9";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"11000b04";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"012a07a9";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"000c07a9";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"0d008d04";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"ff8a07a9";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"000607a9";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"ff7207a9";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"05157930";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"02019c1c";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"09003e0c";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"050a7008";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"08004104";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"002307a9";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"ff8507a9";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"008e07a9";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"14004108";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"08003e04";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"ff9e07a9";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"00b907a9";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"00ff6004";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"002707a9";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"ff8b07a9";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"08003f08";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"1f027704";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"ffcb07a9";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"007f07a9";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"0d008b08";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"0a000104";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"000e07a9";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"ff6507a9";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"002407a9";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"15f71a08";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"07fb6b04";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"007107a9";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"ff8707a9";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"009c07a9";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"0501c328";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"05ffaf14";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"0f005b08";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"0b00d104";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"00460835";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"ff8c0835";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"1f028704";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"ff650835";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"14003104";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"00420835";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"ff7e0835";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"03fe850c";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"08004408";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"01fd3304";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"00e70835";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"fff40835";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"ff9c0835";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"12005404";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"ff730835";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"00170835";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"0519b418";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"020d4d14";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"030bbc10";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"1afb5b08";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"05098504";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"ffa30835";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"003b0835";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"12005304";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"00480835";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"ffd70835";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"ff990835";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"ff930835";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"15f6f904";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"00020835";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"00980835";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"05002d1c";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"0e004d14";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"05ffaf0c";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"1f028704";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"ff6608c9";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"1603b904";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"ff8208c9";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"004b08c9";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"0c006704";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"004408c9";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"ff8d08c9";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"00fd7104";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"004308c9";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"ff8e08c9";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"05157924";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"0a03671c";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"1300880c";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"00fc7f04";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"004a08c9";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"050e1d04";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"ff7008c9";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"ffd608c9";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"10001708";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"05063404";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"fff208c9";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"00a608c9";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"01fc9204";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"003d08c9";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"ffda08c9";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"10033e04";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"00c608c9";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"ffe008c9";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"15f71a08";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"07fb6b04";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"006008c9";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"ff9808c9";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"009308c9";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"05002d1c";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"0f005b08";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"0b00d104";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"00480955";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"ff910955";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"05ffaf0c";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"1f028704";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"ff670955";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"14003104";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"004b0955";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"ff850955";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"0c006704";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"00490955";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"ff930955";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"05157920";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"0a036718";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"03093c10";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"05063408";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"08004604";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"000c0955";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"ff890955";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"0e002204";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"ff990955";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"003b0955";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"14003b04";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"fff70955";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"ff790955";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"10033e04";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"00b40955";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"ffe30955";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"15f71a08";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"18006904";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"ffaf0955";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"00540955";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"008f0955";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"05002d1c";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"0e004d14";
		wait for Clk_period;
		Addr <=  "0001001010111";
		Trees_din <= x"05ffaf0c";
		wait for Clk_period;
		Addr <=  "0001001011000";
		Trees_din <= x"1f028704";
		wait for Clk_period;
		Addr <=  "0001001011001";
		Trees_din <= x"ff670a11";
		wait for Clk_period;
		Addr <=  "0001001011010";
		Trees_din <= x"05fe5404";
		wait for Clk_period;
		Addr <=  "0001001011011";
		Trees_din <= x"ff890a11";
		wait for Clk_period;
		Addr <=  "0001001011100";
		Trees_din <= x"00490a11";
		wait for Clk_period;
		Addr <=  "0001001011101";
		Trees_din <= x"09003904";
		wait for Clk_period;
		Addr <=  "0001001011110";
		Trees_din <= x"00480a11";
		wait for Clk_period;
		Addr <=  "0001001011111";
		Trees_din <= x"ff940a11";
		wait for Clk_period;
		Addr <=  "0001001100000";
		Trees_din <= x"00fd7104";
		wait for Clk_period;
		Addr <=  "0001001100001";
		Trees_din <= x"00480a11";
		wait for Clk_period;
		Addr <=  "0001001100010";
		Trees_din <= x"ff960a11";
		wait for Clk_period;
		Addr <=  "0001001100011";
		Trees_din <= x"0519b43c";
		wait for Clk_period;
		Addr <=  "0001001100100";
		Trees_din <= x"02ffe420";
		wait for Clk_period;
		Addr <=  "0001001100101";
		Trees_din <= x"09003d10";
		wait for Clk_period;
		Addr <=  "0001001100110";
		Trees_din <= x"05089e08";
		wait for Clk_period;
		Addr <=  "0001001100111";
		Trees_din <= x"16040004";
		wait for Clk_period;
		Addr <=  "0001001101000";
		Trees_din <= x"ff870a11";
		wait for Clk_period;
		Addr <=  "0001001101001";
		Trees_din <= x"004a0a11";
		wait for Clk_period;
		Addr <=  "0001001101010";
		Trees_din <= x"02fe7d04";
		wait for Clk_period;
		Addr <=  "0001001101011";
		Trees_din <= x"ffc70a11";
		wait for Clk_period;
		Addr <=  "0001001101100";
		Trees_din <= x"00a10a11";
		wait for Clk_period;
		Addr <=  "0001001101101";
		Trees_din <= x"01fd7808";
		wait for Clk_period;
		Addr <=  "0001001101110";
		Trees_din <= x"03045f04";
		wait for Clk_period;
		Addr <=  "0001001101111";
		Trees_din <= x"00a80a11";
		wait for Clk_period;
		Addr <=  "0001001110000";
		Trees_din <= x"ffd70a11";
		wait for Clk_period;
		Addr <=  "0001001110001";
		Trees_din <= x"14004104";
		wait for Clk_period;
		Addr <=  "0001001110010";
		Trees_din <= x"00510a11";
		wait for Clk_period;
		Addr <=  "0001001110011";
		Trees_din <= x"ffad0a11";
		wait for Clk_period;
		Addr <=  "0001001110100";
		Trees_din <= x"17030d0c";
		wait for Clk_period;
		Addr <=  "0001001110101";
		Trees_din <= x"03054204";
		wait for Clk_period;
		Addr <=  "0001001110110";
		Trees_din <= x"ff960a11";
		wait for Clk_period;
		Addr <=  "0001001110111";
		Trees_din <= x"11006604";
		wait for Clk_period;
		Addr <=  "0001001111000";
		Trees_din <= x"00830a11";
		wait for Clk_period;
		Addr <=  "0001001111001";
		Trees_din <= x"001d0a11";
		wait for Clk_period;
		Addr <=  "0001001111010";
		Trees_din <= x"10010808";
		wait for Clk_period;
		Addr <=  "0001001111011";
		Trees_din <= x"10001904";
		wait for Clk_period;
		Addr <=  "0001001111100";
		Trees_din <= x"fff20a11";
		wait for Clk_period;
		Addr <=  "0001001111101";
		Trees_din <= x"ff730a11";
		wait for Clk_period;
		Addr <=  "0001001111110";
		Trees_din <= x"15f8df04";
		wait for Clk_period;
		Addr <=  "0001001111111";
		Trees_din <= x"00530a11";
		wait for Clk_period;
		Addr <=  "0001010000000";
		Trees_din <= x"ffe30a11";
		wait for Clk_period;
		Addr <=  "0001010000001";
		Trees_din <= x"1c024104";
		wait for Clk_period;
		Addr <=  "0001010000010";
		Trees_din <= x"00180a11";
		wait for Clk_period;
		Addr <=  "0001010000011";
		Trees_din <= x"008c0a11";
		wait for Clk_period;
		Addr <=  "0001010000100";
		Trees_din <= x"05ffaf14";
		wait for Clk_period;
		Addr <=  "0001010000101";
		Trees_din <= x"0f005b08";
		wait for Clk_period;
		Addr <=  "0001010000110";
		Trees_din <= x"15f73704";
		wait for Clk_period;
		Addr <=  "0001010000111";
		Trees_din <= x"ff9e0aad";
		wait for Clk_period;
		Addr <=  "0001010001000";
		Trees_din <= x"004a0aad";
		wait for Clk_period;
		Addr <=  "0001010001001";
		Trees_din <= x"1f028704";
		wait for Clk_period;
		Addr <=  "0001010001010";
		Trees_din <= x"ff680aad";
		wait for Clk_period;
		Addr <=  "0001010001011";
		Trees_din <= x"00fd8504";
		wait for Clk_period;
		Addr <=  "0001010001100";
		Trees_din <= x"004b0aad";
		wait for Clk_period;
		Addr <=  "0001010001101";
		Trees_din <= x"ff8b0aad";
		wait for Clk_period;
		Addr <=  "0001010001110";
		Trees_din <= x"050f8828";
		wait for Clk_period;
		Addr <=  "0001010001111";
		Trees_din <= x"0305bc14";
		wait for Clk_period;
		Addr <=  "0001010010000";
		Trees_din <= x"04044110";
		wait for Clk_period;
		Addr <=  "0001010010001";
		Trees_din <= x"0c006408";
		wait for Clk_period;
		Addr <=  "0001010010010";
		Trees_din <= x"1300b804";
		wait for Clk_period;
		Addr <=  "0001010010011";
		Trees_din <= x"ffac0aad";
		wait for Clk_period;
		Addr <=  "0001010010100";
		Trees_din <= x"00550aad";
		wait for Clk_period;
		Addr <=  "0001010010101";
		Trees_din <= x"1703e304";
		wait for Clk_period;
		Addr <=  "0001010010110";
		Trees_din <= x"00060aad";
		wait for Clk_period;
		Addr <=  "0001010010111";
		Trees_din <= x"00a30aad";
		wait for Clk_period;
		Addr <=  "0001010011000";
		Trees_din <= x"ff860aad";
		wait for Clk_period;
		Addr <=  "0001010011001";
		Trees_din <= x"060c170c";
		wait for Clk_period;
		Addr <=  "0001010011010";
		Trees_din <= x"050e1d08";
		wait for Clk_period;
		Addr <=  "0001010011011";
		Trees_din <= x"01012c04";
		wait for Clk_period;
		Addr <=  "0001010011100";
		Trees_din <= x"ff670aad";
		wait for Clk_period;
		Addr <=  "0001010011101";
		Trees_din <= x"ffed0aad";
		wait for Clk_period;
		Addr <=  "0001010011110";
		Trees_din <= x"fffb0aad";
		wait for Clk_period;
		Addr <=  "0001010011111";
		Trees_din <= x"0507ce04";
		wait for Clk_period;
		Addr <=  "0001010100000";
		Trees_din <= x"ff9d0aad";
		wait for Clk_period;
		Addr <=  "0001010100001";
		Trees_din <= x"00740aad";
		wait for Clk_period;
		Addr <=  "0001010100010";
		Trees_din <= x"15f71d08";
		wait for Clk_period;
		Addr <=  "0001010100011";
		Trees_din <= x"08004b04";
		wait for Clk_period;
		Addr <=  "0001010100100";
		Trees_din <= x"00430aad";
		wait for Clk_period;
		Addr <=  "0001010100101";
		Trees_din <= x"ffb70aad";
		wait for Clk_period;
		Addr <=  "0001010100110";
		Trees_din <= x"0e004408";
		wait for Clk_period;
		Addr <=  "0001010100111";
		Trees_din <= x"0f006f04";
		wait for Clk_period;
		Addr <=  "0001010101000";
		Trees_din <= x"00360aad";
		wait for Clk_period;
		Addr <=  "0001010101001";
		Trees_din <= x"00910aad";
		wait for Clk_period;
		Addr <=  "0001010101010";
		Trees_din <= x"fff30aad";
		wait for Clk_period;
		Addr <=  "0001010101011";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0001010101100";
		Trees_din <= x"05ffaf14";
		wait for Clk_period;
		Addr <=  "0001010101101";
		Trees_din <= x"0f005b08";
		wait for Clk_period;
		Addr <=  "0001010101110";
		Trees_din <= x"12005404";
		wait for Clk_period;
		Addr <=  "0001010101111";
		Trees_din <= x"00490b65";
		wait for Clk_period;
		Addr <=  "0001010110000";
		Trees_din <= x"ffa00b65";
		wait for Clk_period;
		Addr <=  "0001010110001";
		Trees_din <= x"1f028704";
		wait for Clk_period;
		Addr <=  "0001010110010";
		Trees_din <= x"ff690b65";
		wait for Clk_period;
		Addr <=  "0001010110011";
		Trees_din <= x"08003f04";
		wait for Clk_period;
		Addr <=  "0001010110100";
		Trees_din <= x"004c0b65";
		wait for Clk_period;
		Addr <=  "0001010110101";
		Trees_din <= x"ff8e0b65";
		wait for Clk_period;
		Addr <=  "0001010110110";
		Trees_din <= x"0519b440";
		wait for Clk_period;
		Addr <=  "0001010110111";
		Trees_din <= x"0d007020";
		wait for Clk_period;
		Addr <=  "0001010111000";
		Trees_din <= x"01fd9610";
		wait for Clk_period;
		Addr <=  "0001010111001";
		Trees_din <= x"03045f08";
		wait for Clk_period;
		Addr <=  "0001010111010";
		Trees_din <= x"060b0c04";
		wait for Clk_period;
		Addr <=  "0001010111011";
		Trees_din <= x"00b80b65";
		wait for Clk_period;
		Addr <=  "0001010111100";
		Trees_din <= x"000c0b65";
		wait for Clk_period;
		Addr <=  "0001010111101";
		Trees_din <= x"08004404";
		wait for Clk_period;
		Addr <=  "0001010111110";
		Trees_din <= x"ffc10b65";
		wait for Clk_period;
		Addr <=  "0001010111111";
		Trees_din <= x"002a0b65";
		wait for Clk_period;
		Addr <=  "0001011000000";
		Trees_din <= x"0d006e08";
		wait for Clk_period;
		Addr <=  "0001011000001";
		Trees_din <= x"00fc7f04";
		wait for Clk_period;
		Addr <=  "0001011000010";
		Trees_din <= x"00540b65";
		wait for Clk_period;
		Addr <=  "0001011000011";
		Trees_din <= x"ffae0b65";
		wait for Clk_period;
		Addr <=  "0001011000100";
		Trees_din <= x"0505c804";
		wait for Clk_period;
		Addr <=  "0001011000101";
		Trees_din <= x"00180b65";
		wait for Clk_period;
		Addr <=  "0001011000110";
		Trees_din <= x"00860b65";
		wait for Clk_period;
		Addr <=  "0001011000111";
		Trees_din <= x"0505c810";
		wait for Clk_period;
		Addr <=  "0001011001000";
		Trees_din <= x"01fc4e08";
		wait for Clk_period;
		Addr <=  "0001011001001";
		Trees_din <= x"04ffd804";
		wait for Clk_period;
		Addr <=  "0001011001010";
		Trees_din <= x"ff9c0b65";
		wait for Clk_period;
		Addr <=  "0001011001011";
		Trees_din <= x"00740b65";
		wait for Clk_period;
		Addr <=  "0001011001100";
		Trees_din <= x"16021504";
		wait for Clk_period;
		Addr <=  "0001011001101";
		Trees_din <= x"000e0b65";
		wait for Clk_period;
		Addr <=  "0001011001110";
		Trees_din <= x"ff710b65";
		wait for Clk_period;
		Addr <=  "0001011001111";
		Trees_din <= x"1d025a08";
		wait for Clk_period;
		Addr <=  "0001011010000";
		Trees_din <= x"1703f104";
		wait for Clk_period;
		Addr <=  "0001011010001";
		Trees_din <= x"ff780b65";
		wait for Clk_period;
		Addr <=  "0001011010010";
		Trees_din <= x"00090b65";
		wait for Clk_period;
		Addr <=  "0001011010011";
		Trees_din <= x"0c00c804";
		wait for Clk_period;
		Addr <=  "0001011010100";
		Trees_din <= x"ffe50b65";
		wait for Clk_period;
		Addr <=  "0001011010101";
		Trees_din <= x"00520b65";
		wait for Clk_period;
		Addr <=  "0001011010110";
		Trees_din <= x"1d024704";
		wait for Clk_period;
		Addr <=  "0001011010111";
		Trees_din <= x"00170b65";
		wait for Clk_period;
		Addr <=  "0001011011000";
		Trees_din <= x"00840b65";
		wait for Clk_period;
		Addr <=  "0001011011001";
		Trees_din <= x"05ffaf14";
		wait for Clk_period;
		Addr <=  "0001011011010";
		Trees_din <= x"0e004d0c";
		wait for Clk_period;
		Addr <=  "0001011011011";
		Trees_din <= x"00fcc808";
		wait for Clk_period;
		Addr <=  "0001011011100";
		Trees_din <= x"1b027c04";
		wait for Clk_period;
		Addr <=  "0001011011101";
		Trees_din <= x"ff940bf9";
		wait for Clk_period;
		Addr <=  "0001011011110";
		Trees_din <= x"004b0bf9";
		wait for Clk_period;
		Addr <=  "0001011011111";
		Trees_din <= x"ff690bf9";
		wait for Clk_period;
		Addr <=  "0001011100000";
		Trees_din <= x"03fcb204";
		wait for Clk_period;
		Addr <=  "0001011100001";
		Trees_din <= x"004a0bf9";
		wait for Clk_period;
		Addr <=  "0001011100010";
		Trees_din <= x"ffa60bf9";
		wait for Clk_period;
		Addr <=  "0001011100011";
		Trees_din <= x"051d1034";
		wait for Clk_period;
		Addr <=  "0001011100100";
		Trees_din <= x"0d007018";
		wait for Clk_period;
		Addr <=  "0001011100101";
		Trees_din <= x"06ef7508";
		wait for Clk_period;
		Addr <=  "0001011100110";
		Trees_din <= x"0104e104";
		wait for Clk_period;
		Addr <=  "0001011100111";
		Trees_din <= x"ff790bf9";
		wait for Clk_period;
		Addr <=  "0001011101000";
		Trees_din <= x"fffa0bf9";
		wait for Clk_period;
		Addr <=  "0001011101001";
		Trees_din <= x"060c5808";
		wait for Clk_period;
		Addr <=  "0001011101010";
		Trees_din <= x"03093c04";
		wait for Clk_period;
		Addr <=  "0001011101011";
		Trees_din <= x"005b0bf9";
		wait for Clk_period;
		Addr <=  "0001011101100";
		Trees_din <= x"ffbe0bf9";
		wait for Clk_period;
		Addr <=  "0001011101101";
		Trees_din <= x"00fe5004";
		wait for Clk_period;
		Addr <=  "0001011101110";
		Trees_din <= x"ffa50bf9";
		wait for Clk_period;
		Addr <=  "0001011101111";
		Trees_din <= x"fff50bf9";
		wait for Clk_period;
		Addr <=  "0001011110000";
		Trees_din <= x"0506340c";
		wait for Clk_period;
		Addr <=  "0001011110001";
		Trees_din <= x"11001704";
		wait for Clk_period;
		Addr <=  "0001011110010";
		Trees_din <= x"ff750bf9";
		wait for Clk_period;
		Addr <=  "0001011110011";
		Trees_din <= x"15f79004";
		wait for Clk_period;
		Addr <=  "0001011110100";
		Trees_din <= x"008b0bf9";
		wait for Clk_period;
		Addr <=  "0001011110101";
		Trees_din <= x"ffca0bf9";
		wait for Clk_period;
		Addr <=  "0001011110110";
		Trees_din <= x"04fb4b08";
		wait for Clk_period;
		Addr <=  "0001011110111";
		Trees_din <= x"1702b404";
		wait for Clk_period;
		Addr <=  "0001011111000";
		Trees_din <= x"007b0bf9";
		wait for Clk_period;
		Addr <=  "0001011111001";
		Trees_din <= x"ffc80bf9";
		wait for Clk_period;
		Addr <=  "0001011111010";
		Trees_din <= x"1300b504";
		wait for Clk_period;
		Addr <=  "0001011111011";
		Trees_din <= x"ffe30bf9";
		wait for Clk_period;
		Addr <=  "0001011111100";
		Trees_din <= x"00a40bf9";
		wait for Clk_period;
		Addr <=  "0001011111101";
		Trees_din <= x"007f0bf9";
		wait for Clk_period;
		Addr <=  "0001011111110";
		Trees_din <= x"05ffaf14";
		wait for Clk_period;
		Addr <=  "0001011111111";
		Trees_din <= x"0e004d0c";
		wait for Clk_period;
		Addr <=  "0001100000000";
		Trees_din <= x"1f028704";
		wait for Clk_period;
		Addr <=  "0001100000001";
		Trees_din <= x"ff6a0cbd";
		wait for Clk_period;
		Addr <=  "0001100000010";
		Trees_din <= x"09003b04";
		wait for Clk_period;
		Addr <=  "0001100000011";
		Trees_din <= x"00470cbd";
		wait for Clk_period;
		Addr <=  "0001100000100";
		Trees_din <= x"ff9a0cbd";
		wait for Clk_period;
		Addr <=  "0001100000101";
		Trees_din <= x"16040004";
		wait for Clk_period;
		Addr <=  "0001100000110";
		Trees_din <= x"ffa80cbd";
		wait for Clk_period;
		Addr <=  "0001100000111";
		Trees_din <= x"00490cbd";
		wait for Clk_period;
		Addr <=  "0001100001000";
		Trees_din <= x"04f84d24";
		wait for Clk_period;
		Addr <=  "0001100001001";
		Trees_din <= x"1603df0c";
		wait for Clk_period;
		Addr <=  "0001100001010";
		Trees_din <= x"0f006e04";
		wait for Clk_period;
		Addr <=  "0001100001011";
		Trees_din <= x"ffe90cbd";
		wait for Clk_period;
		Addr <=  "0001100001100";
		Trees_din <= x"18004c04";
		wait for Clk_period;
		Addr <=  "0001100001101";
		Trees_din <= x"00180cbd";
		wait for Clk_period;
		Addr <=  "0001100001110";
		Trees_din <= x"00860cbd";
		wait for Clk_period;
		Addr <=  "0001100001111";
		Trees_din <= x"15f7e910";
		wait for Clk_period;
		Addr <=  "0001100010000";
		Trees_din <= x"01ff0f08";
		wait for Clk_period;
		Addr <=  "0001100010001";
		Trees_din <= x"13009a04";
		wait for Clk_period;
		Addr <=  "0001100010010";
		Trees_din <= x"ff9d0cbd";
		wait for Clk_period;
		Addr <=  "0001100010011";
		Trees_din <= x"000f0cbd";
		wait for Clk_period;
		Addr <=  "0001100010100";
		Trees_din <= x"15f6f904";
		wait for Clk_period;
		Addr <=  "0001100010101";
		Trees_din <= x"fff60cbd";
		wait for Clk_period;
		Addr <=  "0001100010110";
		Trees_din <= x"00680cbd";
		wait for Clk_period;
		Addr <=  "0001100010111";
		Trees_din <= x"17037804";
		wait for Clk_period;
		Addr <=  "0001100011000";
		Trees_din <= x"002e0cbd";
		wait for Clk_period;
		Addr <=  "0001100011001";
		Trees_din <= x"ff8c0cbd";
		wait for Clk_period;
		Addr <=  "0001100011010";
		Trees_din <= x"0303d420";
		wait for Clk_period;
		Addr <=  "0001100011011";
		Trees_din <= x"01fd3310";
		wait for Clk_period;
		Addr <=  "0001100011100";
		Trees_din <= x"0e002808";
		wait for Clk_period;
		Addr <=  "0001100011101";
		Trees_din <= x"0e002204";
		wait for Clk_period;
		Addr <=  "0001100011110";
		Trees_din <= x"00490cbd";
		wait for Clk_period;
		Addr <=  "0001100011111";
		Trees_din <= x"ff770cbd";
		wait for Clk_period;
		Addr <=  "0001100100000";
		Trees_din <= x"0b009704";
		wait for Clk_period;
		Addr <=  "0001100100001";
		Trees_din <= x"ffc70cbd";
		wait for Clk_period;
		Addr <=  "0001100100010";
		Trees_din <= x"008a0cbd";
		wait for Clk_period;
		Addr <=  "0001100100011";
		Trees_din <= x"07fed208";
		wait for Clk_period;
		Addr <=  "0001100100100";
		Trees_din <= x"05034004";
		wait for Clk_period;
		Addr <=  "0001100100101";
		Trees_din <= x"ff950cbd";
		wait for Clk_period;
		Addr <=  "0001100100110";
		Trees_din <= x"007c0cbd";
		wait for Clk_period;
		Addr <=  "0001100100111";
		Trees_din <= x"18006804";
		wait for Clk_period;
		Addr <=  "0001100101000";
		Trees_din <= x"00080cbd";
		wait for Clk_period;
		Addr <=  "0001100101001";
		Trees_din <= x"ff720cbd";
		wait for Clk_period;
		Addr <=  "0001100101010";
		Trees_din <= x"07ff1108";
		wait for Clk_period;
		Addr <=  "0001100101011";
		Trees_din <= x"06f8e104";
		wait for Clk_period;
		Addr <=  "0001100101100";
		Trees_din <= x"ffd70cbd";
		wait for Clk_period;
		Addr <=  "0001100101101";
		Trees_din <= x"ff710cbd";
		wait for Clk_period;
		Addr <=  "0001100101110";
		Trees_din <= x"000a0cbd";
		wait for Clk_period;
		Addr <=  "0001100101111";
		Trees_din <= x"05ffaf14";
		wait for Clk_period;
		Addr <=  "0001100110000";
		Trees_din <= x"0f005b08";
		wait for Clk_period;
		Addr <=  "0001100110001";
		Trees_din <= x"03fcb204";
		wait for Clk_period;
		Addr <=  "0001100110010";
		Trees_din <= x"004b0d49";
		wait for Clk_period;
		Addr <=  "0001100110011";
		Trees_din <= x"ffaa0d49";
		wait for Clk_period;
		Addr <=  "0001100110100";
		Trees_din <= x"00fcc808";
		wait for Clk_period;
		Addr <=  "0001100110101";
		Trees_din <= x"1b027c04";
		wait for Clk_period;
		Addr <=  "0001100110110";
		Trees_din <= x"ff9e0d49";
		wait for Clk_period;
		Addr <=  "0001100110111";
		Trees_din <= x"004c0d49";
		wait for Clk_period;
		Addr <=  "0001100111000";
		Trees_din <= x"ff6b0d49";
		wait for Clk_period;
		Addr <=  "0001100111001";
		Trees_din <= x"051d1030";
		wait for Clk_period;
		Addr <=  "0001100111010";
		Trees_din <= x"00ff871c";
		wait for Clk_period;
		Addr <=  "0001100111011";
		Trees_din <= x"1100c010";
		wait for Clk_period;
		Addr <=  "0001100111100";
		Trees_din <= x"0d007108";
		wait for Clk_period;
		Addr <=  "0001100111101";
		Trees_din <= x"060c5804";
		wait for Clk_period;
		Addr <=  "0001100111110";
		Trees_din <= x"005f0d49";
		wait for Clk_period;
		Addr <=  "0001100111111";
		Trees_din <= x"ffce0d49";
		wait for Clk_period;
		Addr <=  "0001101000000";
		Trees_din <= x"14003b04";
		wait for Clk_period;
		Addr <=  "0001101000001";
		Trees_din <= x"001f0d49";
		wait for Clk_period;
		Addr <=  "0001101000010";
		Trees_din <= x"ffae0d49";
		wait for Clk_period;
		Addr <=  "0001101000011";
		Trees_din <= x"1101a604";
		wait for Clk_period;
		Addr <=  "0001101000100";
		Trees_din <= x"ff7e0d49";
		wait for Clk_period;
		Addr <=  "0001101000101";
		Trees_din <= x"0b00d004";
		wait for Clk_period;
		Addr <=  "0001101000110";
		Trees_din <= x"00520d49";
		wait for Clk_period;
		Addr <=  "0001101000111";
		Trees_din <= x"ffe80d49";
		wait for Clk_period;
		Addr <=  "0001101001000";
		Trees_din <= x"0c01e00c";
		wait for Clk_period;
		Addr <=  "0001101001001";
		Trees_din <= x"0d006e04";
		wait for Clk_period;
		Addr <=  "0001101001010";
		Trees_din <= x"ff7c0d49";
		wait for Clk_period;
		Addr <=  "0001101001011";
		Trees_din <= x"01ff9204";
		wait for Clk_period;
		Addr <=  "0001101001100";
		Trees_din <= x"ff9f0d49";
		wait for Clk_period;
		Addr <=  "0001101001101";
		Trees_din <= x"00030d49";
		wait for Clk_period;
		Addr <=  "0001101001110";
		Trees_din <= x"05098504";
		wait for Clk_period;
		Addr <=  "0001101001111";
		Trees_din <= x"ffd00d49";
		wait for Clk_period;
		Addr <=  "0001101010000";
		Trees_din <= x"006f0d49";
		wait for Clk_period;
		Addr <=  "0001101010001";
		Trees_din <= x"00780d49";
		wait for Clk_period;
		Addr <=  "0001101010010";
		Trees_din <= x"05ffaf0c";
		wait for Clk_period;
		Addr <=  "0001101010011";
		Trees_din <= x"060a3604";
		wait for Clk_period;
		Addr <=  "0001101010100";
		Trees_din <= x"ff6c0dcd";
		wait for Clk_period;
		Addr <=  "0001101010101";
		Trees_din <= x"08003f04";
		wait for Clk_period;
		Addr <=  "0001101010110";
		Trees_din <= x"00730dcd";
		wait for Clk_period;
		Addr <=  "0001101010111";
		Trees_din <= x"ff800dcd";
		wait for Clk_period;
		Addr <=  "0001101011000";
		Trees_din <= x"05157930";
		wait for Clk_period;
		Addr <=  "0001101011001";
		Trees_din <= x"02019c20";
		wait for Clk_period;
		Addr <=  "0001101011010";
		Trees_din <= x"050a7010";
		wait for Clk_period;
		Addr <=  "0001101011011";
		Trees_din <= x"0303d408";
		wait for Clk_period;
		Addr <=  "0001101011100";
		Trees_din <= x"0e002704";
		wait for Clk_period;
		Addr <=  "0001101011101";
		Trees_din <= x"ffc20dcd";
		wait for Clk_period;
		Addr <=  "0001101011110";
		Trees_din <= x"00290dcd";
		wait for Clk_period;
		Addr <=  "0001101011111";
		Trees_din <= x"15f76804";
		wait for Clk_period;
		Addr <=  "0001101100000";
		Trees_din <= x"000e0dcd";
		wait for Clk_period;
		Addr <=  "0001101100001";
		Trees_din <= x"ff850dcd";
		wait for Clk_period;
		Addr <=  "0001101100010";
		Trees_din <= x"0d006708";
		wait for Clk_period;
		Addr <=  "0001101100011";
		Trees_din <= x"0b00b804";
		wait for Clk_period;
		Addr <=  "0001101100100";
		Trees_din <= x"ff990dcd";
		wait for Clk_period;
		Addr <=  "0001101100101";
		Trees_din <= x"00360dcd";
		wait for Clk_period;
		Addr <=  "0001101100110";
		Trees_din <= x"0a000904";
		wait for Clk_period;
		Addr <=  "0001101100111";
		Trees_din <= x"00240dcd";
		wait for Clk_period;
		Addr <=  "0001101101000";
		Trees_din <= x"008c0dcd";
		wait for Clk_period;
		Addr <=  "0001101101001";
		Trees_din <= x"0d008c0c";
		wait for Clk_period;
		Addr <=  "0001101101010";
		Trees_din <= x"08003d04";
		wait for Clk_period;
		Addr <=  "0001101101011";
		Trees_din <= x"00130dcd";
		wait for Clk_period;
		Addr <=  "0001101101100";
		Trees_din <= x"1e025404";
		wait for Clk_period;
		Addr <=  "0001101101101";
		Trees_din <= x"ffe40dcd";
		wait for Clk_period;
		Addr <=  "0001101101110";
		Trees_din <= x"ff790dcd";
		wait for Clk_period;
		Addr <=  "0001101101111";
		Trees_din <= x"00310dcd";
		wait for Clk_period;
		Addr <=  "0001101110000";
		Trees_din <= x"15f71a04";
		wait for Clk_period;
		Addr <=  "0001101110001";
		Trees_din <= x"fff30dcd";
		wait for Clk_period;
		Addr <=  "0001101110010";
		Trees_din <= x"00780dcd";
		wait for Clk_period;
		Addr <=  "0001101110011";
		Trees_din <= x"05ffaf0c";
		wait for Clk_period;
		Addr <=  "0001101110100";
		Trees_din <= x"00fd7108";
		wait for Clk_period;
		Addr <=  "0001101110101";
		Trees_din <= x"08003f04";
		wait for Clk_period;
		Addr <=  "0001101110110";
		Trees_din <= x"00940e71";
		wait for Clk_period;
		Addr <=  "0001101110111";
		Trees_din <= x"ff810e71";
		wait for Clk_period;
		Addr <=  "0001101111000";
		Trees_din <= x"ff6d0e71";
		wait for Clk_period;
		Addr <=  "0001101111001";
		Trees_din <= x"04f84d20";
		wait for Clk_period;
		Addr <=  "0001101111010";
		Trees_din <= x"17031a08";
		wait for Clk_period;
		Addr <=  "0001101111011";
		Trees_din <= x"1100ae04";
		wait for Clk_period;
		Addr <=  "0001101111100";
		Trees_din <= x"00840e71";
		wait for Clk_period;
		Addr <=  "0001101111101";
		Trees_din <= x"fff30e71";
		wait for Clk_period;
		Addr <=  "0001101111110";
		Trees_din <= x"1f027c10";
		wait for Clk_period;
		Addr <=  "0001101111111";
		Trees_din <= x"01ff0f08";
		wait for Clk_period;
		Addr <=  "0001110000000";
		Trees_din <= x"19000304";
		wait for Clk_period;
		Addr <=  "0001110000001";
		Trees_din <= x"ffb10e71";
		wait for Clk_period;
		Addr <=  "0001110000010";
		Trees_din <= x"002e0e71";
		wait for Clk_period;
		Addr <=  "0001110000011";
		Trees_din <= x"08003e04";
		wait for Clk_period;
		Addr <=  "0001110000100";
		Trees_din <= x"ffe10e71";
		wait for Clk_period;
		Addr <=  "0001110000101";
		Trees_din <= x"005a0e71";
		wait for Clk_period;
		Addr <=  "0001110000110";
		Trees_din <= x"11006d04";
		wait for Clk_period;
		Addr <=  "0001110000111";
		Trees_din <= x"ff920e71";
		wait for Clk_period;
		Addr <=  "0001110001000";
		Trees_din <= x"fff20e71";
		wait for Clk_period;
		Addr <=  "0001110001001";
		Trees_din <= x"0303d420";
		wait for Clk_period;
		Addr <=  "0001110001010";
		Trees_din <= x"01fd3310";
		wait for Clk_period;
		Addr <=  "0001110001011";
		Trees_din <= x"1300ae08";
		wait for Clk_period;
		Addr <=  "0001110001100";
		Trees_din <= x"0c005f04";
		wait for Clk_period;
		Addr <=  "0001110001101";
		Trees_din <= x"ffa90e71";
		wait for Clk_period;
		Addr <=  "0001110001110";
		Trees_din <= x"00810e71";
		wait for Clk_period;
		Addr <=  "0001110001111";
		Trees_din <= x"0d008004";
		wait for Clk_period;
		Addr <=  "0001110010000";
		Trees_din <= x"ff7a0e71";
		wait for Clk_period;
		Addr <=  "0001110010001";
		Trees_din <= x"00510e71";
		wait for Clk_period;
		Addr <=  "0001110010010";
		Trees_din <= x"03028a08";
		wait for Clk_period;
		Addr <=  "0001110010011";
		Trees_din <= x"06fbc904";
		wait for Clk_period;
		Addr <=  "0001110010100";
		Trees_din <= x"001c0e71";
		wait for Clk_period;
		Addr <=  "0001110010101";
		Trees_din <= x"ff920e71";
		wait for Clk_period;
		Addr <=  "0001110010110";
		Trees_din <= x"07ff4104";
		wait for Clk_period;
		Addr <=  "0001110010111";
		Trees_din <= x"006f0e71";
		wait for Clk_period;
		Addr <=  "0001110011000";
		Trees_din <= x"ffa40e71";
		wait for Clk_period;
		Addr <=  "0001110011001";
		Trees_din <= x"07ff1104";
		wait for Clk_period;
		Addr <=  "0001110011010";
		Trees_din <= x"ff870e71";
		wait for Clk_period;
		Addr <=  "0001110011011";
		Trees_din <= x"000c0e71";
		wait for Clk_period;
		Addr <=  "0001110011100";
		Trees_din <= x"05ffaf0c";
		wait for Clk_period;
		Addr <=  "0001110011101";
		Trees_din <= x"060a3604";
		wait for Clk_period;
		Addr <=  "0001110011110";
		Trees_din <= x"ff6f0f0d";
		wait for Clk_period;
		Addr <=  "0001110011111";
		Trees_din <= x"07ffa904";
		wait for Clk_period;
		Addr <=  "0001110100000";
		Trees_din <= x"ff850f0d";
		wait for Clk_period;
		Addr <=  "0001110100001";
		Trees_din <= x"00820f0d";
		wait for Clk_period;
		Addr <=  "0001110100010";
		Trees_din <= x"05043c1c";
		wait for Clk_period;
		Addr <=  "0001110100011";
		Trees_din <= x"03000310";
		wait for Clk_period;
		Addr <=  "0001110100100";
		Trees_din <= x"01fde40c";
		wait for Clk_period;
		Addr <=  "0001110100101";
		Trees_din <= x"0401c404";
		wait for Clk_period;
		Addr <=  "0001110100110";
		Trees_din <= x"ffe10f0d";
		wait for Clk_period;
		Addr <=  "0001110100111";
		Trees_din <= x"0d006e04";
		wait for Clk_period;
		Addr <=  "0001110101000";
		Trees_din <= x"00900f0d";
		wait for Clk_period;
		Addr <=  "0001110101001";
		Trees_din <= x"fff70f0d";
		wait for Clk_period;
		Addr <=  "0001110101010";
		Trees_din <= x"ff9a0f0d";
		wait for Clk_period;
		Addr <=  "0001110101011";
		Trees_din <= x"1d025108";
		wait for Clk_period;
		Addr <=  "0001110101100";
		Trees_din <= x"05034004";
		wait for Clk_period;
		Addr <=  "0001110101101";
		Trees_din <= x"ffb00f0d";
		wait for Clk_period;
		Addr <=  "0001110101110";
		Trees_din <= x"00550f0d";
		wait for Clk_period;
		Addr <=  "0001110101111";
		Trees_din <= x"ff7c0f0d";
		wait for Clk_period;
		Addr <=  "0001110110000";
		Trees_din <= x"1d02420c";
		wait for Clk_period;
		Addr <=  "0001110110001";
		Trees_din <= x"1602bc04";
		wait for Clk_period;
		Addr <=  "0001110110010";
		Trees_din <= x"001a0f0d";
		wait for Clk_period;
		Addr <=  "0001110110011";
		Trees_din <= x"07fb6b04";
		wait for Clk_period;
		Addr <=  "0001110110100";
		Trees_din <= x"fffa0f0d";
		wait for Clk_period;
		Addr <=  "0001110110101";
		Trees_din <= x"ff930f0d";
		wait for Clk_period;
		Addr <=  "0001110110110";
		Trees_din <= x"1afbe30c";
		wait for Clk_period;
		Addr <=  "0001110110111";
		Trees_din <= x"1603f008";
		wait for Clk_period;
		Addr <=  "0001110111000";
		Trees_din <= x"1100c004";
		wait for Clk_period;
		Addr <=  "0001110111001";
		Trees_din <= x"00510f0d";
		wait for Clk_period;
		Addr <=  "0001110111010";
		Trees_din <= x"ffc50f0d";
		wait for Clk_period;
		Addr <=  "0001110111011";
		Trees_din <= x"ffa30f0d";
		wait for Clk_period;
		Addr <=  "0001110111100";
		Trees_din <= x"09003f08";
		wait for Clk_period;
		Addr <=  "0001110111101";
		Trees_din <= x"10004504";
		wait for Clk_period;
		Addr <=  "0001110111110";
		Trees_din <= x"00410f0d";
		wait for Clk_period;
		Addr <=  "0001110111111";
		Trees_din <= x"ffc80f0d";
		wait for Clk_period;
		Addr <=  "0001111000000";
		Trees_din <= x"14004304";
		wait for Clk_period;
		Addr <=  "0001111000001";
		Trees_din <= x"008f0f0d";
		wait for Clk_period;
		Addr <=  "0001111000010";
		Trees_din <= x"00160f0d";
		wait for Clk_period;
		Addr <=  "0001111000011";
		Trees_din <= x"05ffaf0c";
		wait for Clk_period;
		Addr <=  "0001111000100";
		Trees_din <= x"00fd7108";
		wait for Clk_period;
		Addr <=  "0001111000101";
		Trees_din <= x"01fd4a04";
		wait for Clk_period;
		Addr <=  "0001111000110";
		Trees_din <= x"00950f81";
		wait for Clk_period;
		Addr <=  "0001111000111";
		Trees_din <= x"ff870f81";
		wait for Clk_period;
		Addr <=  "0001111001000";
		Trees_din <= x"ff700f81";
		wait for Clk_period;
		Addr <=  "0001111001001";
		Trees_din <= x"051d102c";
		wait for Clk_period;
		Addr <=  "0001111001010";
		Trees_din <= x"00ff8718";
		wait for Clk_period;
		Addr <=  "0001111001011";
		Trees_din <= x"1100c010";
		wait for Clk_period;
		Addr <=  "0001111001100";
		Trees_din <= x"08004c08";
		wait for Clk_period;
		Addr <=  "0001111001101";
		Trees_din <= x"1300c504";
		wait for Clk_period;
		Addr <=  "0001111001110";
		Trees_din <= x"003e0f81";
		wait for Clk_period;
		Addr <=  "0001111001111";
		Trees_din <= x"ffd60f81";
		wait for Clk_period;
		Addr <=  "0001111010000";
		Trees_din <= x"0b005a04";
		wait for Clk_period;
		Addr <=  "0001111010001";
		Trees_din <= x"00330f81";
		wait for Clk_period;
		Addr <=  "0001111010010";
		Trees_din <= x"ff980f81";
		wait for Clk_period;
		Addr <=  "0001111010011";
		Trees_din <= x"1101a604";
		wait for Clk_period;
		Addr <=  "0001111010100";
		Trees_din <= x"ff8c0f81";
		wait for Clk_period;
		Addr <=  "0001111010101";
		Trees_din <= x"001e0f81";
		wait for Clk_period;
		Addr <=  "0001111010110";
		Trees_din <= x"0c01e00c";
		wait for Clk_period;
		Addr <=  "0001111010111";
		Trees_din <= x"0a000104";
		wait for Clk_period;
		Addr <=  "0001111011000";
		Trees_din <= x"00110f81";
		wait for Clk_period;
		Addr <=  "0001111011001";
		Trees_din <= x"0f007504";
		wait for Clk_period;
		Addr <=  "0001111011010";
		Trees_din <= x"ff820f81";
		wait for Clk_period;
		Addr <=  "0001111011011";
		Trees_din <= x"ffdd0f81";
		wait for Clk_period;
		Addr <=  "0001111011100";
		Trees_din <= x"09003e04";
		wait for Clk_period;
		Addr <=  "0001111011101";
		Trees_din <= x"00420f81";
		wait for Clk_period;
		Addr <=  "0001111011110";
		Trees_din <= x"00090f81";
		wait for Clk_period;
		Addr <=  "0001111011111";
		Trees_din <= x"006c0f81";
		wait for Clk_period;
		Addr <=  "0001111100000";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  4
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"0003ad68";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"00003a34";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"00ff601c";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"1200330c";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"0c002604";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"00ca0125";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"1300dc04";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"00130125";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"ff6b0125";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"00fec408";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"12006304";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"ff520125";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"ffa00125";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"02f88d04";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"00370125";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"ff660125";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"1ffdb408";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"00ffa904";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"ff900125";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"014f0125";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"00ff8f08";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"1002f504";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"ffad0125";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"01090125";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"04049404";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"ff540125";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"ffc00125";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"06ff7b14";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"06f53804";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"ff550125";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"1000d808";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"02f83404";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"00370125";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"ff6e0125";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"1603c304";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"ffbf0125";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"01290125";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"00016510";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"1703ff08";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"03fc6104";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"00420125";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"ff8b0125";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"0f006504";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"ff880125";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"019e0125";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"07047c08";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"06080c04";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"022b0125";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"ff840125";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"02f9d304";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"00ca0125";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"ff790125";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"0501e618";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"0709490c";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"020d4d08";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"1af92904";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"012b0125";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"040b0125";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"ffa40125";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"0009bd08";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"02fa1204";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"00370125";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"ff7c0125";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"02b90125";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"00103e10";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"0503f708";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"01ffb304";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"ff960125";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"01020125";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"18009404";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"ff570125";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"00370125";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"026e0125";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"00016550";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"00ff6028";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"12003310";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"10001e04";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"00c70249";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"07ffd604";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"ff5e0249";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"0a014104";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"ff6f0249";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"004e0249";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"00fec40c";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"12006304";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"ff580249";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"00fe5d04";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"ff7d0249";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"00340249";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"02f88d04";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"003b0249";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"0b011004";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"ff6d0249";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"000a0249";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"07feb014";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"05fcec08";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"1b025804";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"00da0249";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"ff7c0249";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"0000ff04";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"ff590249";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"0303b804";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"009c0249";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"ff820249";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"0407fd10";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"12004408";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"15f75204";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"00800249";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"ff9a0249";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"0e003a04";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"00890249";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"ffa70249";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"ff5c0249";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"0501e630";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"0003f51c";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"06fe9d0c";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"07001f04";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"00c30249";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"09004104";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"ff660249";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"00030249";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"14004008";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"08003d04";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"00170249";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"019c0249";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"03fc4104";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"011d0249";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"ffcb0249";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"04080d10";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"02069308";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"070be104";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"01bf0249";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"005e0249";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"18005f04";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"00c50249";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"ff8d0249";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"ffeb0249";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"00103e10";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"14004f0c";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"02011108";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"0f007e04";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"ff8b0249";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"00bf0249";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"ff5b0249";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"006c0249";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"01a50249";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"00016558";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"00ff6030";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"12003314";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"07ffd604";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"ff63036d";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"1300e508";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"0b00c904";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"ffa1036d";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"0163036d";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"11019904";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"ff6f036d";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"00bc036d";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"00fec40c";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"12006304";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"ff5c036d";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"08005a04";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"ff83036d";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"0045036d";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"02faf508";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"02fabe04";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"ff73036d";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"006e036d";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"0b004b04";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"002d036d";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"ff60036d";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"04019614";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"00ff7d08";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"09004304";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"ff85036d";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"00d6036d";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"15f6eb04";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"fffb036d";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"08003c04";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"ffc3036d";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"ff5d036d";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"0407fd10";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"12003d08";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"15f76804";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"0036036d";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"ff61036d";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"0d007204";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"ffd6036d";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"0072036d";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"ff61036d";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"07fb7f14";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"0009bd0c";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"0d006408";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"18007b04";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"00b3036d";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"ff8b036d";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"ff5e036d";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"030a2d04";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"0147036d";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"ff81036d";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"0007921c";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"06f8410c";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"0c017004";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"ff5b036d";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"0100e304";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"00c4036d";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"ff77036d";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"1af96f08";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"0a00a104";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"ff77036d";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"0027036d";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"11000104";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"0031036d";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"010d036d";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"02fa8a04";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"001e036d";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"020bd304";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"015f036d";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"0054036d";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"0000da64";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"00ff6030";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"12003310";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"07ffd604";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"ff6704d1";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"04063808";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"02fabb04";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"ffcc04d1";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"00fb04d1";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"ff7e04d1";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"00fec410";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"12006308";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"07038a04";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"ff5d04d1";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"ff8504d1";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"00fe5d04";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"ff8b04d1";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"004304d1";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"02faf508";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"02fabe04";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"ff7904d1";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"006204d1";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"03fac704";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"003004d1";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"ff6404d1";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"02fc2318";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"18005b08";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"05fbbf04";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"fff604d1";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"ff6304d1";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"0d006f08";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"00ffbd04";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"003e04d1";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"ff7104d1";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"01fe8f04";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"009d04d1";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"ff7a04d1";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"1d025410";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"05fd9408";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"09003f04";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"ff9804d1";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"019204d1";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"00ff8204";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"003d04d1";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"ff6e04d1";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"03fcaa08";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"02fd7204";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"ff9504d1";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"004404d1";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"ff5d04d1";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"0303d43c";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"0003f520";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"07047c10";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"05ff5308";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"0c005904";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"016904d1";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"007404d1";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"0c021704";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"ff7004d1";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"00a004d1";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"02f9f608";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"17037c04";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"ff8604d1";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"00a704d1";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"08003e04";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"002d04d1";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"ff6204d1";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"070a2310";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"10005808";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"04037904";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"00ed04d1";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"000d04d1";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"01fbf904";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"fff404d1";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"012504d1";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"0009bd08";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"0407ad04";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"ff8504d1";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"003c04d1";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"00b604d1";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"00103e10";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"0d005b04";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"004904d1";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"02011108";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"07fe9804";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"ff8004d1";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"009104d1";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"ff6004d1";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"00f204d1";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"00003a58";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"00feee20";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"12002c08";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"1b028704";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"ff7c060d";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"00d7060d";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"12006310";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"12003308";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"14002d04";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"ff6a060d";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"0048060d";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"07038a04";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"ff61060d";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"ff8a060d";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"10002d04";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"ff8e060d";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"0040060d";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"0b00db20";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"0b005c10";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"04065608";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"1f024604";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"003f060d";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"ff7b060d";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"04072504";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"0202060d";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"ffa4060d";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"16040008";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"0c01db04";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"ff5e060d";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"ffae060d";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"11000004";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"ff76060d";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"0116060d";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"09004410";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"01fd8c08";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"02fb0004";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"00b2060d";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"ffaf060d";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"1b022a04";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"003b060d";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"ff6f060d";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"19000004";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"01d3060d";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"0034060d";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"0501e634";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"00031a1c";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"0701a110";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"06082608";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"0303b804";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"00da060d";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"ff88060d";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"08003d04";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"00c1060d";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"ff66060d";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"1afb1904";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"ff60060d";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"06020d04";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"ffc3060d";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"0050060d";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"04080d10";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"02069308";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"1300a704";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"009b060d";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"00f7060d";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"11001604";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"ff7b060d";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"0099060d";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"03fbe404";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"ff9c060d";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"002c060d";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"00087204";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"ff63060d";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"050c850c";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"09003804";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"ffff060d";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"15f88a04";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"013e060d";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"0023060d";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"ff83060d";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"00003a5c";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"00feee2c";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"12003314";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"1b028608";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"14002e04";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"ff6b0721";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"003c0721";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"05fdf908";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"08004004";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"00db0721";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"00370721";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"ff9a0721";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"12006310";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"07038a08";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"00fec404";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"ff610721";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"ff8b0721";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"16040004";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"ff6b0721";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"00c20721";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"1c027404";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"ff930721";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"00440721";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"02fc2320";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"0b00db10";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"09004708";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"16040004";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"ff610721";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"00090721";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"1002f504";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"ffd00721";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"01020721";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"09004308";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"11000704";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"00a10721";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"ffb10721";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"02faf804";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"00250721";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"01cc0721";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"03fb2d04";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"00440721";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"19009508";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"06fbc904";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"ffda0721";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"ff6b0721";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"002c0721";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"05089e28";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"00036a14";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"06097710";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"0701a108";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"05ff5304";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"00a90721";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"ffac0721";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"05fb9c04";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"ff680721";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"00040721";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"ff6d0721";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"0213ee10";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"07072708";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"08004f04";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"00d50721";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"00590721";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"0009bd04";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"fff30721";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"00be0721";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"ff940721";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"00103e04";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"ff690721";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"00710721";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"00ff6044";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"12003314";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"07ffd604";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"ff72080d";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"0406380c";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"ffa2080d";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"0a025604";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"011c080d";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"ffaa080d";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"ff90080d";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"00fec418";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"12006310";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"07038a08";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"1f028704";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"ff61080d";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"ff9e080d";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"01fcaf04";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"00c4080d";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"ff6f080d";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"13006b04";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"ff9d080d";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"0044080d";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"02faf50c";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"04050808";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"0d007404";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"00e6080d";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"ff84080d";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"ff69080d";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"09004f08";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"18005a04";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"ffb9080d";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"ff65080d";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"003b080d";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"00079220";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"0303d418";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"060a9910";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"04080d08";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"0f006704";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"ff9a080d";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"004a080d";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"02fe0404";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"ff7b080d";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"001b080d";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"16018204";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"003e080d";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"ff6a080d";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"08003c04";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"ffe6080d";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"ff64080d";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"030a2d10";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"070a2308";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"05089e04";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"00cd080d";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"003d080d";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"04027404";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"008e080d";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"ffa3080d";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"ff8c080d";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"00ff603c";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"00fe7318";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"1cf7ed04";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"001a0915";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"01fbc908";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"0b00ce04";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"ff990915";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"00470915";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"1f028704";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"ff640915";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"1b028704";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"004a0915";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"ff800915";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"08003a08";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"02fad504";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"00f80915";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"ffff0915";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"07ff7e0c";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"02fa9f08";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"1603e004";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"00480915";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"ff900915";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"ff660915";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"02fabe08";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"10030a04";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"ff680915";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"003c0915";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"03fbaf04";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"005f0915";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"ffb20915";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"00031a28";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"04006014";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"0c02520c";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"05fcf504";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"ffdb0915";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"19000704";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"ff630915";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"ffb60915";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"08003f04";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"00a70915";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"ff950915";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"05fb6508";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"00024004";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"ff650915";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"fffa0915";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"060aff08";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"01fe8f04";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"003b0915";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"ffc30915";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"ff760915";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"050c851c";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"06f9a110";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"00066308";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"11013e04";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"ff840915";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"005b0915";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"0009bd04";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"003b0915";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"00ac0915";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"0b00ed08";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"12003504";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"00210915";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"00c70915";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"fffd0915";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"ff7e0915";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"00ff6040";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"00fe731c";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"1cf7ed04";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"001c0a49";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"01fbc908";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"07fece04";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"ff9e0a49";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"00490a49";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"1f028708";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"18004404";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"ffa80a49";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"ff640a49";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"1b028704";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"00460a49";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"ff850a49";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"08003a08";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"0c012a04";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"fffb0a49";
		wait for Clk_period;
		Addr <=  "0001001010111";
		Trees_din <= x"00d10a49";
		wait for Clk_period;
		Addr <=  "0001001011000";
		Trees_din <= x"07ff7e0c";
		wait for Clk_period;
		Addr <=  "0001001011001";
		Trees_din <= x"02fa9f08";
		wait for Clk_period;
		Addr <=  "0001001011010";
		Trees_din <= x"12004304";
		wait for Clk_period;
		Addr <=  "0001001011011";
		Trees_din <= x"00490a49";
		wait for Clk_period;
		Addr <=  "0001001011100";
		Trees_din <= x"ff960a49";
		wait for Clk_period;
		Addr <=  "0001001011101";
		Trees_din <= x"ff690a49";
		wait for Clk_period;
		Addr <=  "0001001011110";
		Trees_din <= x"02fabe08";
		wait for Clk_period;
		Addr <=  "0001001011111";
		Trees_din <= x"10030a04";
		wait for Clk_period;
		Addr <=  "0001001100000";
		Trees_din <= x"ff6b0a49";
		wait for Clk_period;
		Addr <=  "0001001100001";
		Trees_din <= x"00390a49";
		wait for Clk_period;
		Addr <=  "0001001100010";
		Trees_din <= x"02fad204";
		wait for Clk_period;
		Addr <=  "0001001100011";
		Trees_din <= x"00a70a49";
		wait for Clk_period;
		Addr <=  "0001001100100";
		Trees_din <= x"ffc70a49";
		wait for Clk_period;
		Addr <=  "0001001100101";
		Trees_din <= x"00016534";
		wait for Clk_period;
		Addr <=  "0001001100110";
		Trees_din <= x"0f007a1c";
		wait for Clk_period;
		Addr <=  "0001001100111";
		Trees_din <= x"0f00690c";
		wait for Clk_period;
		Addr <=  "0001001101000";
		Trees_din <= x"06096c04";
		wait for Clk_period;
		Addr <=  "0001001101001";
		Trees_din <= x"ff6a0a49";
		wait for Clk_period;
		Addr <=  "0001001101010";
		Trees_din <= x"07fef604";
		wait for Clk_period;
		Addr <=  "0001001101011";
		Trees_din <= x"ffa20a49";
		wait for Clk_period;
		Addr <=  "0001001101100";
		Trees_din <= x"00470a49";
		wait for Clk_period;
		Addr <=  "0001001101101";
		Trees_din <= x"0e003608";
		wait for Clk_period;
		Addr <=  "0001001101110";
		Trees_din <= x"1d027d04";
		wait for Clk_period;
		Addr <=  "0001001101111";
		Trees_din <= x"009d0a49";
		wait for Clk_period;
		Addr <=  "0001001110000";
		Trees_din <= x"ffa30a49";
		wait for Clk_period;
		Addr <=  "0001001110001";
		Trees_din <= x"0f006e04";
		wait for Clk_period;
		Addr <=  "0001001110010";
		Trees_din <= x"00880a49";
		wait for Clk_period;
		Addr <=  "0001001110011";
		Trees_din <= x"ff920a49";
		wait for Clk_period;
		Addr <=  "0001001110100";
		Trees_din <= x"1e028710";
		wait for Clk_period;
		Addr <=  "0001001110101";
		Trees_din <= x"08004a08";
		wait for Clk_period;
		Addr <=  "0001001110110";
		Trees_din <= x"14003004";
		wait for Clk_period;
		Addr <=  "0001001110111";
		Trees_din <= x"ffd10a49";
		wait for Clk_period;
		Addr <=  "0001001111000";
		Trees_din <= x"ff5e0a49";
		wait for Clk_period;
		Addr <=  "0001001111001";
		Trees_din <= x"0e003104";
		wait for Clk_period;
		Addr <=  "0001001111010";
		Trees_din <= x"ffa60a49";
		wait for Clk_period;
		Addr <=  "0001001111011";
		Trees_din <= x"00580a49";
		wait for Clk_period;
		Addr <=  "0001001111100";
		Trees_din <= x"09004004";
		wait for Clk_period;
		Addr <=  "0001001111101";
		Trees_din <= x"ffa40a49";
		wait for Clk_period;
		Addr <=  "0001001111110";
		Trees_din <= x"01150a49";
		wait for Clk_period;
		Addr <=  "0001001111111";
		Trees_din <= x"05089e20";
		wait for Clk_period;
		Addr <=  "0001010000000";
		Trees_din <= x"00079210";
		wait for Clk_period;
		Addr <=  "0001010000001";
		Trees_din <= x"06f84108";
		wait for Clk_period;
		Addr <=  "0001010000010";
		Trees_din <= x"0c017004";
		wait for Clk_period;
		Addr <=  "0001010000011";
		Trees_din <= x"ff660a49";
		wait for Clk_period;
		Addr <=  "0001010000100";
		Trees_din <= x"003e0a49";
		wait for Clk_period;
		Addr <=  "0001010000101";
		Trees_din <= x"12004204";
		wait for Clk_period;
		Addr <=  "0001010000110";
		Trees_din <= x"009b0a49";
		wait for Clk_period;
		Addr <=  "0001010000111";
		Trees_din <= x"00320a49";
		wait for Clk_period;
		Addr <=  "0001010001000";
		Trees_din <= x"070a2308";
		wait for Clk_period;
		Addr <=  "0001010001001";
		Trees_din <= x"1afe7804";
		wait for Clk_period;
		Addr <=  "0001010001010";
		Trees_din <= x"00b50a49";
		wait for Clk_period;
		Addr <=  "0001010001011";
		Trees_din <= x"002a0a49";
		wait for Clk_period;
		Addr <=  "0001010001100";
		Trees_din <= x"04027404";
		wait for Clk_period;
		Addr <=  "0001010001101";
		Trees_din <= x"00730a49";
		wait for Clk_period;
		Addr <=  "0001010001110";
		Trees_din <= x"ffa80a49";
		wait for Clk_period;
		Addr <=  "0001010001111";
		Trees_din <= x"00103e04";
		wait for Clk_period;
		Addr <=  "0001010010000";
		Trees_din <= x"ff760a49";
		wait for Clk_period;
		Addr <=  "0001010010001";
		Trees_din <= x"00550a49";
		wait for Clk_period;
		Addr <=  "0001010010010";
		Trees_din <= x"00ff4740";
		wait for Clk_period;
		Addr <=  "0001010010011";
		Trees_din <= x"00fe731c";
		wait for Clk_period;
		Addr <=  "0001010010100";
		Trees_din <= x"1cf7ed04";
		wait for Clk_period;
		Addr <=  "0001010010101";
		Trees_din <= x"001a0b65";
		wait for Clk_period;
		Addr <=  "0001010010110";
		Trees_din <= x"01fbc908";
		wait for Clk_period;
		Addr <=  "0001010010111";
		Trees_din <= x"08004204";
		wait for Clk_period;
		Addr <=  "0001010011000";
		Trees_din <= x"00470b65";
		wait for Clk_period;
		Addr <=  "0001010011001";
		Trees_din <= x"ffa20b65";
		wait for Clk_period;
		Addr <=  "0001010011010";
		Trees_din <= x"1f028708";
		wait for Clk_period;
		Addr <=  "0001010011011";
		Trees_din <= x"18004404";
		wait for Clk_period;
		Addr <=  "0001010011100";
		Trees_din <= x"ffb00b65";
		wait for Clk_period;
		Addr <=  "0001010011101";
		Trees_din <= x"ff650b65";
		wait for Clk_period;
		Addr <=  "0001010011110";
		Trees_din <= x"1c028704";
		wait for Clk_period;
		Addr <=  "0001010011111";
		Trees_din <= x"00470b65";
		wait for Clk_period;
		Addr <=  "0001010100000";
		Trees_din <= x"ff890b65";
		wait for Clk_period;
		Addr <=  "0001010100001";
		Trees_din <= x"07ff7e0c";
		wait for Clk_period;
		Addr <=  "0001010100010";
		Trees_din <= x"02fa9f08";
		wait for Clk_period;
		Addr <=  "0001010100011";
		Trees_din <= x"07fe9804";
		wait for Clk_period;
		Addr <=  "0001010100100";
		Trees_din <= x"00490b65";
		wait for Clk_period;
		Addr <=  "0001010100101";
		Trees_din <= x"ffa20b65";
		wait for Clk_period;
		Addr <=  "0001010100110";
		Trees_din <= x"ff6b0b65";
		wait for Clk_period;
		Addr <=  "0001010100111";
		Trees_din <= x"08003a08";
		wait for Clk_period;
		Addr <=  "0001010101000";
		Trees_din <= x"16032a04";
		wait for Clk_period;
		Addr <=  "0001010101001";
		Trees_din <= x"00cf0b65";
		wait for Clk_period;
		Addr <=  "0001010101010";
		Trees_din <= x"00060b65";
		wait for Clk_period;
		Addr <=  "0001010101011";
		Trees_din <= x"02fabe08";
		wait for Clk_period;
		Addr <=  "0001010101100";
		Trees_din <= x"10030a04";
		wait for Clk_period;
		Addr <=  "0001010101101";
		Trees_din <= x"ff6e0b65";
		wait for Clk_period;
		Addr <=  "0001010101110";
		Trees_din <= x"00310b65";
		wait for Clk_period;
		Addr <=  "0001010101111";
		Trees_din <= x"02fb0b04";
		wait for Clk_period;
		Addr <=  "0001010110000";
		Trees_din <= x"005a0b65";
		wait for Clk_period;
		Addr <=  "0001010110001";
		Trees_din <= x"ffae0b65";
		wait for Clk_period;
		Addr <=  "0001010110010";
		Trees_din <= x"0001652c";
		wait for Clk_period;
		Addr <=  "0001010110011";
		Trees_din <= x"02fbee18";
		wait for Clk_period;
		Addr <=  "0001010110100";
		Trees_din <= x"04074210";
		wait for Clk_period;
		Addr <=  "0001010110101";
		Trees_din <= x"18005d08";
		wait for Clk_period;
		Addr <=  "0001010110110";
		Trees_din <= x"0f007704";
		wait for Clk_period;
		Addr <=  "0001010110111";
		Trees_din <= x"00980b65";
		wait for Clk_period;
		Addr <=  "0001010111000";
		Trees_din <= x"ff980b65";
		wait for Clk_period;
		Addr <=  "0001010111001";
		Trees_din <= x"17040004";
		wait for Clk_period;
		Addr <=  "0001010111010";
		Trees_din <= x"005d0b65";
		wait for Clk_period;
		Addr <=  "0001010111011";
		Trees_din <= x"ff750b65";
		wait for Clk_period;
		Addr <=  "0001010111100";
		Trees_din <= x"1afa6704";
		wait for Clk_period;
		Addr <=  "0001010111101";
		Trees_din <= x"003b0b65";
		wait for Clk_period;
		Addr <=  "0001010111110";
		Trees_din <= x"ff720b65";
		wait for Clk_period;
		Addr <=  "0001010111111";
		Trees_din <= x"1b027710";
		wait for Clk_period;
		Addr <=  "0001011000000";
		Trees_din <= x"04035808";
		wait for Clk_period;
		Addr <=  "0001011000001";
		Trees_din <= x"04018304";
		wait for Clk_period;
		Addr <=  "0001011000010";
		Trees_din <= x"ffa80b65";
		wait for Clk_period;
		Addr <=  "0001011000011";
		Trees_din <= x"00be0b65";
		wait for Clk_period;
		Addr <=  "0001011000100";
		Trees_din <= x"09004504";
		wait for Clk_period;
		Addr <=  "0001011000101";
		Trees_din <= x"ff6a0b65";
		wait for Clk_period;
		Addr <=  "0001011000110";
		Trees_din <= x"002b0b65";
		wait for Clk_period;
		Addr <=  "0001011000111";
		Trees_din <= x"ff640b65";
		wait for Clk_period;
		Addr <=  "0001011001000";
		Trees_din <= x"05089e1c";
		wait for Clk_period;
		Addr <=  "0001011001001";
		Trees_din <= x"00079210";
		wait for Clk_period;
		Addr <=  "0001011001010";
		Trees_din <= x"0500a708";
		wait for Clk_period;
		Addr <=  "0001011001011";
		Trees_din <= x"12004204";
		wait for Clk_period;
		Addr <=  "0001011001100";
		Trees_din <= x"00820b65";
		wait for Clk_period;
		Addr <=  "0001011001101";
		Trees_din <= x"001e0b65";
		wait for Clk_period;
		Addr <=  "0001011001110";
		Trees_din <= x"09004404";
		wait for Clk_period;
		Addr <=  "0001011001111";
		Trees_din <= x"ff7c0b65";
		wait for Clk_period;
		Addr <=  "0001011010000";
		Trees_din <= x"ffec0b65";
		wait for Clk_period;
		Addr <=  "0001011010001";
		Trees_din <= x"070a2308";
		wait for Clk_period;
		Addr <=  "0001011010010";
		Trees_din <= x"1afe7804";
		wait for Clk_period;
		Addr <=  "0001011010011";
		Trees_din <= x"00aa0b65";
		wait for Clk_period;
		Addr <=  "0001011010100";
		Trees_din <= x"00260b65";
		wait for Clk_period;
		Addr <=  "0001011010101";
		Trees_din <= x"00170b65";
		wait for Clk_period;
		Addr <=  "0001011010110";
		Trees_din <= x"00103e04";
		wait for Clk_period;
		Addr <=  "0001011010111";
		Trees_din <= x"ff7b0b65";
		wait for Clk_period;
		Addr <=  "0001011011000";
		Trees_din <= x"004a0b65";
		wait for Clk_period;
		Addr <=  "0001011011001";
		Trees_din <= x"00feee2c";
		wait for Clk_period;
		Addr <=  "0001011011010";
		Trees_din <= x"12003310";
		wait for Clk_period;
		Addr <=  "0001011011011";
		Trees_din <= x"17032208";
		wait for Clk_period;
		Addr <=  "0001011011100";
		Trees_din <= x"1702be04";
		wait for Clk_period;
		Addr <=  "0001011011101";
		Trees_din <= x"ffa40c41";
		wait for Clk_period;
		Addr <=  "0001011011110";
		Trees_din <= x"00c40c41";
		wait for Clk_period;
		Addr <=  "0001011011111";
		Trees_din <= x"0f009d04";
		wait for Clk_period;
		Addr <=  "0001011100000";
		Trees_din <= x"ff790c41";
		wait for Clk_period;
		Addr <=  "0001011100001";
		Trees_din <= x"00300c41";
		wait for Clk_period;
		Addr <=  "0001011100010";
		Trees_din <= x"12006318";
		wait for Clk_period;
		Addr <=  "0001011100011";
		Trees_din <= x"07038a10";
		wait for Clk_period;
		Addr <=  "0001011100100";
		Trees_din <= x"00fec408";
		wait for Clk_period;
		Addr <=  "0001011100101";
		Trees_din <= x"1f028704";
		wait for Clk_period;
		Addr <=  "0001011100110";
		Trees_din <= x"ff650c41";
		wait for Clk_period;
		Addr <=  "0001011100111";
		Trees_din <= x"ffc00c41";
		wait for Clk_period;
		Addr <=  "0001011101000";
		Trees_din <= x"01fe8504";
		wait for Clk_period;
		Addr <=  "0001011101001";
		Trees_din <= x"ff750c41";
		wait for Clk_period;
		Addr <=  "0001011101010";
		Trees_din <= x"00740c41";
		wait for Clk_period;
		Addr <=  "0001011101011";
		Trees_din <= x"01fcaf04";
		wait for Clk_period;
		Addr <=  "0001011101100";
		Trees_din <= x"00e20c41";
		wait for Clk_period;
		Addr <=  "0001011101101";
		Trees_din <= x"ff7d0c41";
		wait for Clk_period;
		Addr <=  "0001011101110";
		Trees_din <= x"000f0c41";
		wait for Clk_period;
		Addr <=  "0001011101111";
		Trees_din <= x"0003f52c";
		wait for Clk_period;
		Addr <=  "0001011110000";
		Trees_din <= x"04009714";
		wait for Clk_period;
		Addr <=  "0001011110001";
		Trees_din <= x"08003f08";
		wait for Clk_period;
		Addr <=  "0001011110010";
		Trees_din <= x"0c025204";
		wait for Clk_period;
		Addr <=  "0001011110011";
		Trees_din <= x"ff8d0c41";
		wait for Clk_period;
		Addr <=  "0001011110100";
		Trees_din <= x"00a50c41";
		wait for Clk_period;
		Addr <=  "0001011110101";
		Trees_din <= x"0b00f104";
		wait for Clk_period;
		Addr <=  "0001011110110";
		Trees_din <= x"ff660c41";
		wait for Clk_period;
		Addr <=  "0001011110111";
		Trees_din <= x"13009604";
		wait for Clk_period;
		Addr <=  "0001011111000";
		Trees_din <= x"ff9d0c41";
		wait for Clk_period;
		Addr <=  "0001011111001";
		Trees_din <= x"006f0c41";
		wait for Clk_period;
		Addr <=  "0001011111010";
		Trees_din <= x"1300dc10";
		wait for Clk_period;
		Addr <=  "0001011111011";
		Trees_din <= x"0c022008";
		wait for Clk_period;
		Addr <=  "0001011111100";
		Trees_din <= x"01fe8f04";
		wait for Clk_period;
		Addr <=  "0001011111101";
		Trees_din <= x"003b0c41";
		wait for Clk_period;
		Addr <=  "0001011111110";
		Trees_din <= x"ffc00c41";
		wait for Clk_period;
		Addr <=  "0001011111111";
		Trees_din <= x"00014e04";
		wait for Clk_period;
		Addr <=  "0001100000000";
		Trees_din <= x"ff910c41";
		wait for Clk_period;
		Addr <=  "0001100000001";
		Trees_din <= x"003a0c41";
		wait for Clk_period;
		Addr <=  "0001100000010";
		Trees_din <= x"0f00a504";
		wait for Clk_period;
		Addr <=  "0001100000011";
		Trees_din <= x"ff6b0c41";
		wait for Clk_period;
		Addr <=  "0001100000100";
		Trees_din <= x"fff80c41";
		wait for Clk_period;
		Addr <=  "0001100000101";
		Trees_din <= x"050c8514";
		wait for Clk_period;
		Addr <=  "0001100000110";
		Trees_din <= x"0213ee10";
		wait for Clk_period;
		Addr <=  "0001100000111";
		Trees_din <= x"07072708";
		wait for Clk_period;
		Addr <=  "0001100001000";
		Trees_din <= x"09003804";
		wait for Clk_period;
		Addr <=  "0001100001001";
		Trees_din <= x"00340c41";
		wait for Clk_period;
		Addr <=  "0001100001010";
		Trees_din <= x"009d0c41";
		wait for Clk_period;
		Addr <=  "0001100001011";
		Trees_din <= x"01ffbf04";
		wait for Clk_period;
		Addr <=  "0001100001100";
		Trees_din <= x"005a0c41";
		wait for Clk_period;
		Addr <=  "0001100001101";
		Trees_din <= x"ffcb0c41";
		wait for Clk_period;
		Addr <=  "0001100001110";
		Trees_din <= x"ffab0c41";
		wait for Clk_period;
		Addr <=  "0001100001111";
		Trees_din <= x"ff970c41";
		wait for Clk_period;
		Addr <=  "0001100010000";
		Trees_din <= x"00feee24";
		wait for Clk_period;
		Addr <=  "0001100010001";
		Trees_din <= x"1800470c";
		wait for Clk_period;
		Addr <=  "0001100010010";
		Trees_din <= x"14002d08";
		wait for Clk_period;
		Addr <=  "0001100010011";
		Trees_din <= x"1b028804";
		wait for Clk_period;
		Addr <=  "0001100010100";
		Trees_din <= x"ff770ce5";
		wait for Clk_period;
		Addr <=  "0001100010101";
		Trees_din <= x"00710ce5";
		wait for Clk_period;
		Addr <=  "0001100010110";
		Trees_din <= x"00b50ce5";
		wait for Clk_period;
		Addr <=  "0001100010111";
		Trees_din <= x"00fe3604";
		wait for Clk_period;
		Addr <=  "0001100011000";
		Trees_din <= x"ff660ce5";
		wait for Clk_period;
		Addr <=  "0001100011001";
		Trees_din <= x"01fc4508";
		wait for Clk_period;
		Addr <=  "0001100011010";
		Trees_din <= x"10001e04";
		wait for Clk_period;
		Addr <=  "0001100011011";
		Trees_din <= x"00e00ce5";
		wait for Clk_period;
		Addr <=  "0001100011100";
		Trees_din <= x"ffa30ce5";
		wait for Clk_period;
		Addr <=  "0001100011101";
		Trees_din <= x"0a00a104";
		wait for Clk_period;
		Addr <=  "0001100011110";
		Trees_din <= x"ff6b0ce5";
		wait for Clk_period;
		Addr <=  "0001100011111";
		Trees_din <= x"0a016004";
		wait for Clk_period;
		Addr <=  "0001100100000";
		Trees_din <= x"00300ce5";
		wait for Clk_period;
		Addr <=  "0001100100001";
		Trees_din <= x"ff790ce5";
		wait for Clk_period;
		Addr <=  "0001100100010";
		Trees_din <= x"060aff2c";
		wait for Clk_period;
		Addr <=  "0001100100011";
		Trees_din <= x"00079218";
		wait for Clk_period;
		Addr <=  "0001100100100";
		Trees_din <= x"0303d410";
		wait for Clk_period;
		Addr <=  "0001100100101";
		Trees_din <= x"04080d08";
		wait for Clk_period;
		Addr <=  "0001100100110";
		Trees_din <= x"1300dc04";
		wait for Clk_period;
		Addr <=  "0001100100111";
		Trees_din <= x"00270ce5";
		wait for Clk_period;
		Addr <=  "0001100101000";
		Trees_din <= x"ffa20ce5";
		wait for Clk_period;
		Addr <=  "0001100101001";
		Trees_din <= x"15f7b104";
		wait for Clk_period;
		Addr <=  "0001100101010";
		Trees_din <= x"00030ce5";
		wait for Clk_period;
		Addr <=  "0001100101011";
		Trees_din <= x"ff6e0ce5";
		wait for Clk_period;
		Addr <=  "0001100101100";
		Trees_din <= x"08003c04";
		wait for Clk_period;
		Addr <=  "0001100101101";
		Trees_din <= x"fff80ce5";
		wait for Clk_period;
		Addr <=  "0001100101110";
		Trees_din <= x"ff6f0ce5";
		wait for Clk_period;
		Addr <=  "0001100101111";
		Trees_din <= x"0213ee10";
		wait for Clk_period;
		Addr <=  "0001100110000";
		Trees_din <= x"04036d08";
		wait for Clk_period;
		Addr <=  "0001100110001";
		Trees_din <= x"05089e04";
		wait for Clk_period;
		Addr <=  "0001100110010";
		Trees_din <= x"00a50ce5";
		wait for Clk_period;
		Addr <=  "0001100110011";
		Trees_din <= x"00070ce5";
		wait for Clk_period;
		Addr <=  "0001100110100";
		Trees_din <= x"07081904";
		wait for Clk_period;
		Addr <=  "0001100110101";
		Trees_din <= x"006f0ce5";
		wait for Clk_period;
		Addr <=  "0001100110110";
		Trees_din <= x"ffc70ce5";
		wait for Clk_period;
		Addr <=  "0001100110111";
		Trees_din <= x"ffae0ce5";
		wait for Clk_period;
		Addr <=  "0001100111000";
		Trees_din <= x"ff720ce5";
		wait for Clk_period;
		Addr <=  "0001100111001";
		Trees_din <= x"00feee28";
		wait for Clk_period;
		Addr <=  "0001100111010";
		Trees_din <= x"1800470c";
		wait for Clk_period;
		Addr <=  "0001100111011";
		Trees_din <= x"14002d08";
		wait for Clk_period;
		Addr <=  "0001100111100";
		Trees_din <= x"1b028804";
		wait for Clk_period;
		Addr <=  "0001100111101";
		Trees_din <= x"ff7b0dd9";
		wait for Clk_period;
		Addr <=  "0001100111110";
		Trees_din <= x"00650dd9";
		wait for Clk_period;
		Addr <=  "0001100111111";
		Trees_din <= x"00a00dd9";
		wait for Clk_period;
		Addr <=  "0001101000000";
		Trees_din <= x"00fe3604";
		wait for Clk_period;
		Addr <=  "0001101000001";
		Trees_din <= x"ff670dd9";
		wait for Clk_period;
		Addr <=  "0001101000010";
		Trees_din <= x"07038a10";
		wait for Clk_period;
		Addr <=  "0001101000011";
		Trees_din <= x"1f027c08";
		wait for Clk_period;
		Addr <=  "0001101000100";
		Trees_din <= x"0b008d04";
		wait for Clk_period;
		Addr <=  "0001101000101";
		Trees_din <= x"ffe30dd9";
		wait for Clk_period;
		Addr <=  "0001101000110";
		Trees_din <= x"ff6c0dd9";
		wait for Clk_period;
		Addr <=  "0001101000111";
		Trees_din <= x"07008704";
		wait for Clk_period;
		Addr <=  "0001101001000";
		Trees_din <= x"ff830dd9";
		wait for Clk_period;
		Addr <=  "0001101001001";
		Trees_din <= x"007f0dd9";
		wait for Clk_period;
		Addr <=  "0001101001010";
		Trees_din <= x"1703f304";
		wait for Clk_period;
		Addr <=  "0001101001011";
		Trees_din <= x"ffa30dd9";
		wait for Clk_period;
		Addr <=  "0001101001100";
		Trees_din <= x"00df0dd9";
		wait for Clk_period;
		Addr <=  "0001101001101";
		Trees_din <= x"00016520";
		wait for Clk_period;
		Addr <=  "0001101001110";
		Trees_din <= x"14004818";
		wait for Clk_period;
		Addr <=  "0001101001111";
		Trees_din <= x"1400470c";
		wait for Clk_period;
		Addr <=  "0001101010000";
		Trees_din <= x"02f9df04";
		wait for Clk_period;
		Addr <=  "0001101010001";
		Trees_din <= x"ff6a0dd9";
		wait for Clk_period;
		Addr <=  "0001101010010";
		Trees_din <= x"03fc6104";
		wait for Clk_period;
		Addr <=  "0001101010011";
		Trees_din <= x"00440dd9";
		wait for Clk_period;
		Addr <=  "0001101010100";
		Trees_din <= x"ffdf0dd9";
		wait for Clk_period;
		Addr <=  "0001101010101";
		Trees_din <= x"1c027b08";
		wait for Clk_period;
		Addr <=  "0001101010110";
		Trees_din <= x"13008404";
		wait for Clk_period;
		Addr <=  "0001101010111";
		Trees_din <= x"00020dd9";
		wait for Clk_period;
		Addr <=  "0001101011000";
		Trees_din <= x"011c0dd9";
		wait for Clk_period;
		Addr <=  "0001101011001";
		Trees_din <= x"fff10dd9";
		wait for Clk_period;
		Addr <=  "0001101011010";
		Trees_din <= x"07052104";
		wait for Clk_period;
		Addr <=  "0001101011011";
		Trees_din <= x"ff6a0dd9";
		wait for Clk_period;
		Addr <=  "0001101011100";
		Trees_din <= x"00940dd9";
		wait for Clk_period;
		Addr <=  "0001101011101";
		Trees_din <= x"09004720";
		wait for Clk_period;
		Addr <=  "0001101011110";
		Trees_din <= x"09003f10";
		wait for Clk_period;
		Addr <=  "0001101011111";
		Trees_din <= x"05fd4908";
		wait for Clk_period;
		Addr <=  "0001101100000";
		Trees_din <= x"05fcc704";
		wait for Clk_period;
		Addr <=  "0001101100001";
		Trees_din <= x"00200dd9";
		wait for Clk_period;
		Addr <=  "0001101100010";
		Trees_din <= x"00a90dd9";
		wait for Clk_period;
		Addr <=  "0001101100011";
		Trees_din <= x"000d0b04";
		wait for Clk_period;
		Addr <=  "0001101100100";
		Trees_din <= x"ffbf0dd9";
		wait for Clk_period;
		Addr <=  "0001101100101";
		Trees_din <= x"00840dd9";
		wait for Clk_period;
		Addr <=  "0001101100110";
		Trees_din <= x"06023608";
		wait for Clk_period;
		Addr <=  "0001101100111";
		Trees_din <= x"00031a04";
		wait for Clk_period;
		Addr <=  "0001101101000";
		Trees_din <= x"ffdd0dd9";
		wait for Clk_period;
		Addr <=  "0001101101001";
		Trees_din <= x"00760dd9";
		wait for Clk_period;
		Addr <=  "0001101101010";
		Trees_din <= x"14004904";
		wait for Clk_period;
		Addr <=  "0001101101011";
		Trees_din <= x"00da0dd9";
		wait for Clk_period;
		Addr <=  "0001101101100";
		Trees_din <= x"00260dd9";
		wait for Clk_period;
		Addr <=  "0001101101101";
		Trees_din <= x"1001190c";
		wait for Clk_period;
		Addr <=  "0001101101110";
		Trees_din <= x"12004904";
		wait for Clk_period;
		Addr <=  "0001101101111";
		Trees_din <= x"fff30dd9";
		wait for Clk_period;
		Addr <=  "0001101110000";
		Trees_din <= x"0a000904";
		wait for Clk_period;
		Addr <=  "0001101110001";
		Trees_din <= x"ffde0dd9";
		wait for Clk_period;
		Addr <=  "0001101110010";
		Trees_din <= x"ff560dd9";
		wait for Clk_period;
		Addr <=  "0001101110011";
		Trees_din <= x"08004904";
		wait for Clk_period;
		Addr <=  "0001101110100";
		Trees_din <= x"ffd20dd9";
		wait for Clk_period;
		Addr <=  "0001101110101";
		Trees_din <= x"00850dd9";
		wait for Clk_period;
		Addr <=  "0001101110110";
		Trees_din <= x"00feee28";
		wait for Clk_period;
		Addr <=  "0001101110111";
		Trees_din <= x"12003310";
		wait for Clk_period;
		Addr <=  "0001101111000";
		Trees_din <= x"07008e08";
		wait for Clk_period;
		Addr <=  "0001101111001";
		Trees_din <= x"14002d04";
		wait for Clk_period;
		Addr <=  "0001101111010";
		Trees_din <= x"ff870ead";
		wait for Clk_period;
		Addr <=  "0001101111011";
		Trees_din <= x"00210ead";
		wait for Clk_period;
		Addr <=  "0001101111100";
		Trees_din <= x"1b028704";
		wait for Clk_period;
		Addr <=  "0001101111101";
		Trees_din <= x"ffff0ead";
		wait for Clk_period;
		Addr <=  "0001101111110";
		Trees_din <= x"009d0ead";
		wait for Clk_period;
		Addr <=  "0001101111111";
		Trees_din <= x"00fe3604";
		wait for Clk_period;
		Addr <=  "0001110000000";
		Trees_din <= x"ff680ead";
		wait for Clk_period;
		Addr <=  "0001110000001";
		Trees_din <= x"01fc4508";
		wait for Clk_period;
		Addr <=  "0001110000010";
		Trees_din <= x"16040004";
		wait for Clk_period;
		Addr <=  "0001110000011";
		Trees_din <= x"ffa70ead";
		wait for Clk_period;
		Addr <=  "0001110000100";
		Trees_din <= x"00dd0ead";
		wait for Clk_period;
		Addr <=  "0001110000101";
		Trees_din <= x"0a00a104";
		wait for Clk_period;
		Addr <=  "0001110000110";
		Trees_din <= x"ff6e0ead";
		wait for Clk_period;
		Addr <=  "0001110000111";
		Trees_din <= x"06085504";
		wait for Clk_period;
		Addr <=  "0001110001000";
		Trees_din <= x"ff7d0ead";
		wait for Clk_period;
		Addr <=  "0001110001001";
		Trees_din <= x"00480ead";
		wait for Clk_period;
		Addr <=  "0001110001010";
		Trees_din <= x"060aff40";
		wait for Clk_period;
		Addr <=  "0001110001011";
		Trees_din <= x"0b00be20";
		wait for Clk_period;
		Addr <=  "0001110001100";
		Trees_din <= x"03fe5810";
		wait for Clk_period;
		Addr <=  "0001110001101";
		Trees_din <= x"18005f08";
		wait for Clk_period;
		Addr <=  "0001110001110";
		Trees_din <= x"03fcb204";
		wait for Clk_period;
		Addr <=  "0001110001111";
		Trees_din <= x"ff630ead";
		wait for Clk_period;
		Addr <=  "0001110010000";
		Trees_din <= x"fff30ead";
		wait for Clk_period;
		Addr <=  "0001110010001";
		Trees_din <= x"0d007204";
		wait for Clk_period;
		Addr <=  "0001110010010";
		Trees_din <= x"ffce0ead";
		wait for Clk_period;
		Addr <=  "0001110010011";
		Trees_din <= x"00550ead";
		wait for Clk_period;
		Addr <=  "0001110010100";
		Trees_din <= x"00044308";
		wait for Clk_period;
		Addr <=  "0001110010101";
		Trees_din <= x"01fbc904";
		wait for Clk_period;
		Addr <=  "0001110010110";
		Trees_din <= x"002d0ead";
		wait for Clk_period;
		Addr <=  "0001110010111";
		Trees_din <= x"ff7f0ead";
		wait for Clk_period;
		Addr <=  "0001110011000";
		Trees_din <= x"06f6aa04";
		wait for Clk_period;
		Addr <=  "0001110011001";
		Trees_din <= x"ffdf0ead";
		wait for Clk_period;
		Addr <=  "0001110011010";
		Trees_din <= x"00810ead";
		wait for Clk_period;
		Addr <=  "0001110011011";
		Trees_din <= x"0405fc10";
		wait for Clk_period;
		Addr <=  "0001110011100";
		Trees_din <= x"09003c08";
		wait for Clk_period;
		Addr <=  "0001110011101";
		Trees_din <= x"08004104";
		wait for Clk_period;
		Addr <=  "0001110011110";
		Trees_din <= x"ffbd0ead";
		wait for Clk_period;
		Addr <=  "0001110011111";
		Trees_din <= x"003a0ead";
		wait for Clk_period;
		Addr <=  "0001110100000";
		Trees_din <= x"1c026904";
		wait for Clk_period;
		Addr <=  "0001110100001";
		Trees_din <= x"00240ead";
		wait for Clk_period;
		Addr <=  "0001110100010";
		Trees_din <= x"00a50ead";
		wait for Clk_period;
		Addr <=  "0001110100011";
		Trees_din <= x"12003708";
		wait for Clk_period;
		Addr <=  "0001110100100";
		Trees_din <= x"03fcc104";
		wait for Clk_period;
		Addr <=  "0001110100101";
		Trees_din <= x"001a0ead";
		wait for Clk_period;
		Addr <=  "0001110100110";
		Trees_din <= x"00c90ead";
		wait for Clk_period;
		Addr <=  "0001110100111";
		Trees_din <= x"08004304";
		wait for Clk_period;
		Addr <=  "0001110101000";
		Trees_din <= x"ff7c0ead";
		wait for Clk_period;
		Addr <=  "0001110101001";
		Trees_din <= x"002d0ead";
		wait for Clk_period;
		Addr <=  "0001110101010";
		Trees_din <= x"ff770ead";
		wait for Clk_period;
		Addr <=  "0001110101011";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0001110101100";
		Trees_din <= x"00feee2c";
		wait for Clk_period;
		Addr <=  "0001110101101";
		Trees_din <= x"07008710";
		wait for Clk_period;
		Addr <=  "0001110101110";
		Trees_din <= x"00fed508";
		wait for Clk_period;
		Addr <=  "0001110101111";
		Trees_din <= x"08003a04";
		wait for Clk_period;
		Addr <=  "0001110110000";
		Trees_din <= x"ffe90f5d";
		wait for Clk_period;
		Addr <=  "0001110110001";
		Trees_din <= x"ff690f5d";
		wait for Clk_period;
		Addr <=  "0001110110010";
		Trees_din <= x"0b00b904";
		wait for Clk_period;
		Addr <=  "0001110110011";
		Trees_din <= x"004a0f5d";
		wait for Clk_period;
		Addr <=  "0001110110100";
		Trees_din <= x"ffa80f5d";
		wait for Clk_period;
		Addr <=  "0001110110101";
		Trees_din <= x"0700a308";
		wait for Clk_period;
		Addr <=  "0001110110110";
		Trees_din <= x"17032204";
		wait for Clk_period;
		Addr <=  "0001110110111";
		Trees_din <= x"014c0f5d";
		wait for Clk_period;
		Addr <=  "0001110111000";
		Trees_din <= x"ffb00f5d";
		wait for Clk_period;
		Addr <=  "0001110111001";
		Trees_din <= x"01fc4508";
		wait for Clk_period;
		Addr <=  "0001110111010";
		Trees_din <= x"08004204";
		wait for Clk_period;
		Addr <=  "0001110111011";
		Trees_din <= x"00d90f5d";
		wait for Clk_period;
		Addr <=  "0001110111100";
		Trees_din <= x"000e0f5d";
		wait for Clk_period;
		Addr <=  "0001110111101";
		Trees_din <= x"0d009204";
		wait for Clk_period;
		Addr <=  "0001110111110";
		Trees_din <= x"ff6c0f5d";
		wait for Clk_period;
		Addr <=  "0001110111111";
		Trees_din <= x"0d009704";
		wait for Clk_period;
		Addr <=  "0001111000000";
		Trees_din <= x"00990f5d";
		wait for Clk_period;
		Addr <=  "0001111000001";
		Trees_din <= x"ff980f5d";
		wait for Clk_period;
		Addr <=  "0001111000010";
		Trees_din <= x"060aff28";
		wait for Clk_period;
		Addr <=  "0001111000011";
		Trees_din <= x"00079218";
		wait for Clk_period;
		Addr <=  "0001111000100";
		Trees_din <= x"0303d410";
		wait for Clk_period;
		Addr <=  "0001111000101";
		Trees_din <= x"07011008";
		wait for Clk_period;
		Addr <=  "0001111000110";
		Trees_din <= x"1d027604";
		wait for Clk_period;
		Addr <=  "0001111000111";
		Trees_din <= x"005a0f5d";
		wait for Clk_period;
		Addr <=  "0001111001000";
		Trees_din <= x"ffe50f5d";
		wait for Clk_period;
		Addr <=  "0001111001001";
		Trees_din <= x"01ffcd04";
		wait for Clk_period;
		Addr <=  "0001111001010";
		Trees_din <= x"00000f5d";
		wait for Clk_period;
		Addr <=  "0001111001011";
		Trees_din <= x"ff760f5d";
		wait for Clk_period;
		Addr <=  "0001111001100";
		Trees_din <= x"0b00ed04";
		wait for Clk_period;
		Addr <=  "0001111001101";
		Trees_din <= x"ff750f5d";
		wait for Clk_period;
		Addr <=  "0001111001110";
		Trees_din <= x"ffe50f5d";
		wait for Clk_period;
		Addr <=  "0001111001111";
		Trees_din <= x"0107cc0c";
		wait for Clk_period;
		Addr <=  "0001111010000";
		Trees_din <= x"0402a804";
		wait for Clk_period;
		Addr <=  "0001111010001";
		Trees_din <= x"008b0f5d";
		wait for Clk_period;
		Addr <=  "0001111010010";
		Trees_din <= x"07081904";
		wait for Clk_period;
		Addr <=  "0001111010011";
		Trees_din <= x"006e0f5d";
		wait for Clk_period;
		Addr <=  "0001111010100";
		Trees_din <= x"ffc10f5d";
		wait for Clk_period;
		Addr <=  "0001111010101";
		Trees_din <= x"fffb0f5d";
		wait for Clk_period;
		Addr <=  "0001111010110";
		Trees_din <= x"ff7b0f5d";
		wait for Clk_period;
		Addr <=  "0001111010111";
		Trees_din <= x"00feee2c";
		wait for Clk_period;
		Addr <=  "0001111011000";
		Trees_din <= x"07008710";
		wait for Clk_period;
		Addr <=  "0001111011001";
		Trees_din <= x"00fed508";
		wait for Clk_period;
		Addr <=  "0001111011010";
		Trees_din <= x"08003a04";
		wait for Clk_period;
		Addr <=  "0001111011011";
		Trees_din <= x"ffec1061";
		wait for Clk_period;
		Addr <=  "0001111011100";
		Trees_din <= x"ff691061";
		wait for Clk_period;
		Addr <=  "0001111011101";
		Trees_din <= x"1300b104";
		wait for Clk_period;
		Addr <=  "0001111011110";
		Trees_din <= x"ffaa1061";
		wait for Clk_period;
		Addr <=  "0001111011111";
		Trees_din <= x"00491061";
		wait for Clk_period;
		Addr <=  "0001111100000";
		Trees_din <= x"0700a308";
		wait for Clk_period;
		Addr <=  "0001111100001";
		Trees_din <= x"08004204";
		wait for Clk_period;
		Addr <=  "0001111100010";
		Trees_din <= x"01221061";
		wait for Clk_period;
		Addr <=  "0001111100011";
		Trees_din <= x"ffb01061";
		wait for Clk_period;
		Addr <=  "0001111100100";
		Trees_din <= x"01fc4508";
		wait for Clk_period;
		Addr <=  "0001111100101";
		Trees_din <= x"10000b04";
		wait for Clk_period;
		Addr <=  "0001111100110";
		Trees_din <= x"00ed1061";
		wait for Clk_period;
		Addr <=  "0001111100111";
		Trees_din <= x"ffb11061";
		wait for Clk_period;
		Addr <=  "0001111101000";
		Trees_din <= x"0d009204";
		wait for Clk_period;
		Addr <=  "0001111101001";
		Trees_din <= x"ff6e1061";
		wait for Clk_period;
		Addr <=  "0001111101010";
		Trees_din <= x"0d009704";
		wait for Clk_period;
		Addr <=  "0001111101011";
		Trees_din <= x"00881061";
		wait for Clk_period;
		Addr <=  "0001111101100";
		Trees_din <= x"ff9d1061";
		wait for Clk_period;
		Addr <=  "0001111101101";
		Trees_din <= x"00016524";
		wait for Clk_period;
		Addr <=  "0001111101110";
		Trees_din <= x"0407fd20";
		wait for Clk_period;
		Addr <=  "0001111101111";
		Trees_din <= x"03fc6110";
		wait for Clk_period;
		Addr <=  "0001111110000";
		Trees_din <= x"11000208";
		wait for Clk_period;
		Addr <=  "0001111110001";
		Trees_din <= x"10006604";
		wait for Clk_period;
		Addr <=  "0001111110010";
		Trees_din <= x"ff721061";
		wait for Clk_period;
		Addr <=  "0001111110011";
		Trees_din <= x"00271061";
		wait for Clk_period;
		Addr <=  "0001111110100";
		Trees_din <= x"16040004";
		wait for Clk_period;
		Addr <=  "0001111110101";
		Trees_din <= x"00261061";
		wait for Clk_period;
		Addr <=  "0001111110110";
		Trees_din <= x"01211061";
		wait for Clk_period;
		Addr <=  "0001111110111";
		Trees_din <= x"1b027508";
		wait for Clk_period;
		Addr <=  "0001111111000";
		Trees_din <= x"1e027004";
		wait for Clk_period;
		Addr <=  "0001111111001";
		Trees_din <= x"ffe51061";
		wait for Clk_period;
		Addr <=  "0001111111010";
		Trees_din <= x"00731061";
		wait for Clk_period;
		Addr <=  "0001111111011";
		Trees_din <= x"00ff0c04";
		wait for Clk_period;
		Addr <=  "0001111111100";
		Trees_din <= x"006d1061";
		wait for Clk_period;
		Addr <=  "0001111111101";
		Trees_din <= x"ff821061";
		wait for Clk_period;
		Addr <=  "0001111111110";
		Trees_din <= x"ff771061";
		wait for Clk_period;
		Addr <=  "0001111111111";
		Trees_din <= x"10009c1c";
		wait for Clk_period;
		Addr <=  "0010000000000";
		Trees_din <= x"0a002310";
		wait for Clk_period;
		Addr <=  "0010000000001";
		Trees_din <= x"0b00c408";
		wait for Clk_period;
		Addr <=  "0010000000010";
		Trees_din <= x"06fb6604";
		wait for Clk_period;
		Addr <=  "0010000000011";
		Trees_din <= x"fff51061";
		wait for Clk_period;
		Addr <=  "0010000000100";
		Trees_din <= x"00d51061";
		wait for Clk_period;
		Addr <=  "0010000000101";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "0010000000110";
		Trees_din <= x"006e1061";
		wait for Clk_period;
		Addr <=  "0010000000111";
		Trees_din <= x"ffd71061";
		wait for Clk_period;
		Addr <=  "0010000001000";
		Trees_din <= x"11001e08";
		wait for Clk_period;
		Addr <=  "0010000001001";
		Trees_din <= x"0405f104";
		wait for Clk_period;
		Addr <=  "0010000001010";
		Trees_din <= x"00231061";
		wait for Clk_period;
		Addr <=  "0010000001011";
		Trees_din <= x"ff781061";
		wait for Clk_period;
		Addr <=  "0010000001100";
		Trees_din <= x"ff501061";
		wait for Clk_period;
		Addr <=  "0010000001101";
		Trees_din <= x"0300950c";
		wait for Clk_period;
		Addr <=  "0010000001110";
		Trees_din <= x"07021904";
		wait for Clk_period;
		Addr <=  "0010000001111";
		Trees_din <= x"00c51061";
		wait for Clk_period;
		Addr <=  "0010000010000";
		Trees_din <= x"1300a204";
		wait for Clk_period;
		Addr <=  "0010000010001";
		Trees_din <= x"ffbb1061";
		wait for Clk_period;
		Addr <=  "0010000010010";
		Trees_din <= x"00641061";
		wait for Clk_period;
		Addr <=  "0010000010011";
		Trees_din <= x"09004708";
		wait for Clk_period;
		Addr <=  "0010000010100";
		Trees_din <= x"11001104";
		wait for Clk_period;
		Addr <=  "0010000010101";
		Trees_din <= x"006c1061";
		wait for Clk_period;
		Addr <=  "0010000010110";
		Trees_din <= x"ffe31061";
		wait for Clk_period;
		Addr <=  "0010000010111";
		Trees_din <= x"ff821061";
		wait for Clk_period;
		Addr <=  "0010000011000";
		Trees_din <= x"00feee30";
		wait for Clk_period;
		Addr <=  "0010000011001";
		Trees_din <= x"00fe360c";
		wait for Clk_period;
		Addr <=  "0010000011010";
		Trees_din <= x"18004408";
		wait for Clk_period;
		Addr <=  "0010000011011";
		Trees_din <= x"07008104";
		wait for Clk_period;
		Addr <=  "0010000011100";
		Trees_din <= x"ffa31165";
		wait for Clk_period;
		Addr <=  "0010000011101";
		Trees_din <= x"00681165";
		wait for Clk_period;
		Addr <=  "0010000011110";
		Trees_din <= x"ff6b1165";
		wait for Clk_period;
		Addr <=  "0010000011111";
		Trees_din <= x"08004118";
		wait for Clk_period;
		Addr <=  "0010000100000";
		Trees_din <= x"07008708";
		wait for Clk_period;
		Addr <=  "0010000100001";
		Trees_din <= x"19001504";
		wait for Clk_period;
		Addr <=  "0010000100010";
		Trees_din <= x"ff891165";
		wait for Clk_period;
		Addr <=  "0010000100011";
		Trees_din <= x"00221165";
		wait for Clk_period;
		Addr <=  "0010000100100";
		Trees_din <= x"08003f08";
		wait for Clk_period;
		Addr <=  "0010000100101";
		Trees_din <= x"1d028404";
		wait for Clk_period;
		Addr <=  "0010000100110";
		Trees_din <= x"ffa61165";
		wait for Clk_period;
		Addr <=  "0010000100111";
		Trees_din <= x"00181165";
		wait for Clk_period;
		Addr <=  "0010000101000";
		Trees_din <= x"05fdd804";
		wait for Clk_period;
		Addr <=  "0010000101001";
		Trees_din <= x"00211165";
		wait for Clk_period;
		Addr <=  "0010000101010";
		Trees_din <= x"01641165";
		wait for Clk_period;
		Addr <=  "0010000101011";
		Trees_din <= x"12004f04";
		wait for Clk_period;
		Addr <=  "0010000101100";
		Trees_din <= x"ff731165";
		wait for Clk_period;
		Addr <=  "0010000101101";
		Trees_din <= x"14004704";
		wait for Clk_period;
		Addr <=  "0010000101110";
		Trees_din <= x"00b11165";
		wait for Clk_period;
		Addr <=  "0010000101111";
		Trees_din <= x"ff911165";
		wait for Clk_period;
		Addr <=  "0010000110000";
		Trees_din <= x"0003f530";
		wait for Clk_period;
		Addr <=  "0010000110001";
		Trees_din <= x"04006010";
		wait for Clk_period;
		Addr <=  "0010000110010";
		Trees_din <= x"08003f08";
		wait for Clk_period;
		Addr <=  "0010000110011";
		Trees_din <= x"0c025204";
		wait for Clk_period;
		Addr <=  "0010000110100";
		Trees_din <= x"ffa11165";
		wait for Clk_period;
		Addr <=  "0010000110101";
		Trees_din <= x"00871165";
		wait for Clk_period;
		Addr <=  "0010000110110";
		Trees_din <= x"0b00f104";
		wait for Clk_period;
		Addr <=  "0010000110111";
		Trees_din <= x"ff6e1165";
		wait for Clk_period;
		Addr <=  "0010000111000";
		Trees_din <= x"ffd51165";
		wait for Clk_period;
		Addr <=  "0010000111001";
		Trees_din <= x"0c023a10";
		wait for Clk_period;
		Addr <=  "0010000111010";
		Trees_din <= x"0f006708";
		wait for Clk_period;
		Addr <=  "0010000111011";
		Trees_din <= x"0f005704";
		wait for Clk_period;
		Addr <=  "0010000111100";
		Trees_din <= x"00531165";
		wait for Clk_period;
		Addr <=  "0010000111101";
		Trees_din <= x"ff6b1165";
		wait for Clk_period;
		Addr <=  "0010000111110";
		Trees_din <= x"1300dc04";
		wait for Clk_period;
		Addr <=  "0010000111111";
		Trees_din <= x"00281165";
		wait for Clk_period;
		Addr <=  "0010001000000";
		Trees_din <= x"ff911165";
		wait for Clk_period;
		Addr <=  "0010001000001";
		Trees_din <= x"0000ee08";
		wait for Clk_period;
		Addr <=  "0010001000010";
		Trees_din <= x"0f008604";
		wait for Clk_period;
		Addr <=  "0010001000011";
		Trees_din <= x"ff691165";
		wait for Clk_period;
		Addr <=  "0010001000100";
		Trees_din <= x"001e1165";
		wait for Clk_period;
		Addr <=  "0010001000101";
		Trees_din <= x"0d006904";
		wait for Clk_period;
		Addr <=  "0010001000110";
		Trees_din <= x"00881165";
		wait for Clk_period;
		Addr <=  "0010001000111";
		Trees_din <= x"ff991165";
		wait for Clk_period;
		Addr <=  "0010001001000";
		Trees_din <= x"02069314";
		wait for Clk_period;
		Addr <=  "0010001001001";
		Trees_din <= x"19000b0c";
		wait for Clk_period;
		Addr <=  "0010001001010";
		Trees_din <= x"01fea604";
		wait for Clk_period;
		Addr <=  "0010001001011";
		Trees_din <= x"00941165";
		wait for Clk_period;
		Addr <=  "0010001001100";
		Trees_din <= x"0009bd04";
		wait for Clk_period;
		Addr <=  "0010001001101";
		Trees_din <= x"ffea1165";
		wait for Clk_period;
		Addr <=  "0010001001110";
		Trees_din <= x"007e1165";
		wait for Clk_period;
		Addr <=  "0010001001111";
		Trees_din <= x"01fdc804";
		wait for Clk_period;
		Addr <=  "0010001010000";
		Trees_din <= x"ffb01165";
		wait for Clk_period;
		Addr <=  "0010001010001";
		Trees_din <= x"004c1165";
		wait for Clk_period;
		Addr <=  "0010001010010";
		Trees_din <= x"00087208";
		wait for Clk_period;
		Addr <=  "0010001010011";
		Trees_din <= x"020bd304";
		wait for Clk_period;
		Addr <=  "0010001010100";
		Trees_din <= x"ff921165";
		wait for Clk_period;
		Addr <=  "0010001010101";
		Trees_din <= x"fff41165";
		wait for Clk_period;
		Addr <=  "0010001010110";
		Trees_din <= x"14004604";
		wait for Clk_period;
		Addr <=  "0010001010111";
		Trees_din <= x"ffeb1165";
		wait for Clk_period;
		Addr <=  "0010001011000";
		Trees_din <= x"00561165";
		wait for Clk_period;
		Addr <=  "0010001011001";
		Trees_din <= x"00fe360c";
		wait for Clk_period;
		Addr <=  "0010001011010";
		Trees_din <= x"18004408";
		wait for Clk_period;
		Addr <=  "0010001011011";
		Trees_din <= x"07008104";
		wait for Clk_period;
		Addr <=  "0010001011100";
		Trees_din <= x"ffa711e9";
		wait for Clk_period;
		Addr <=  "0010001011101";
		Trees_din <= x"005d11e9";
		wait for Clk_period;
		Addr <=  "0010001011110";
		Trees_din <= x"ff6c11e9";
		wait for Clk_period;
		Addr <=  "0010001011111";
		Trees_din <= x"060aff34";
		wait for Clk_period;
		Addr <=  "0010001100000";
		Trees_din <= x"04058320";
		wait for Clk_period;
		Addr <=  "0010001100001";
		Trees_din <= x"0b00ba10";
		wait for Clk_period;
		Addr <=  "0010001100010";
		Trees_din <= x"0404a808";
		wait for Clk_period;
		Addr <=  "0010001100011";
		Trees_din <= x"10001704";
		wait for Clk_period;
		Addr <=  "0010001100100";
		Trees_din <= x"002911e9";
		wait for Clk_period;
		Addr <=  "0010001100101";
		Trees_din <= x"ffaf11e9";
		wait for Clk_period;
		Addr <=  "0010001100110";
		Trees_din <= x"05fdbe04";
		wait for Clk_period;
		Addr <=  "0010001100111";
		Trees_din <= x"009b11e9";
		wait for Clk_period;
		Addr <=  "0010001101000";
		Trees_din <= x"ff7f11e9";
		wait for Clk_period;
		Addr <=  "0010001101001";
		Trees_din <= x"05ff5308";
		wait for Clk_period;
		Addr <=  "0010001101010";
		Trees_din <= x"08004704";
		wait for Clk_period;
		Addr <=  "0010001101011";
		Trees_din <= x"005511e9";
		wait for Clk_period;
		Addr <=  "0010001101100";
		Trees_din <= x"ffc911e9";
		wait for Clk_period;
		Addr <=  "0010001101101";
		Trees_din <= x"0c017f04";
		wait for Clk_period;
		Addr <=  "0010001101110";
		Trees_din <= x"ff9a11e9";
		wait for Clk_period;
		Addr <=  "0010001101111";
		Trees_din <= x"003411e9";
		wait for Clk_period;
		Addr <=  "0010001110000";
		Trees_din <= x"09004f10";
		wait for Clk_period;
		Addr <=  "0010001110001";
		Trees_din <= x"00fff308";
		wait for Clk_period;
		Addr <=  "0010001110010";
		Trees_din <= x"0d006004";
		wait for Clk_period;
		Addr <=  "0010001110011";
		Trees_din <= x"003c11e9";
		wait for Clk_period;
		Addr <=  "0010001110100";
		Trees_din <= x"ff8011e9";
		wait for Clk_period;
		Addr <=  "0010001110101";
		Trees_din <= x"10009a04";
		wait for Clk_period;
		Addr <=  "0010001110110";
		Trees_din <= x"ffd211e9";
		wait for Clk_period;
		Addr <=  "0010001110111";
		Trees_din <= x"004a11e9";
		wait for Clk_period;
		Addr <=  "0010001111000";
		Trees_din <= x"00d311e9";
		wait for Clk_period;
		Addr <=  "0010001111001";
		Trees_din <= x"ff7711e9";
		wait for Clk_period;
		Addr <=  "0010001111010";
		Trees_din <= x"00fe360c";
		wait for Clk_period;
		Addr <=  "0010001111011";
		Trees_din <= x"18004408";
		wait for Clk_period;
		Addr <=  "0010001111100";
		Trees_din <= x"07008104";
		wait for Clk_period;
		Addr <=  "0010001111101";
		Trees_din <= x"ffab1245";
		wait for Clk_period;
		Addr <=  "0010001111110";
		Trees_din <= x"00561245";
		wait for Clk_period;
		Addr <=  "0010001111111";
		Trees_din <= x"ff6d1245";
		wait for Clk_period;
		Addr <=  "0010010000000";
		Trees_din <= x"060aff20";
		wait for Clk_period;
		Addr <=  "0010010000001";
		Trees_din <= x"0009bd18";
		wait for Clk_period;
		Addr <=  "0010010000010";
		Trees_din <= x"0303d410";
		wait for Clk_period;
		Addr <=  "0010010000011";
		Trees_din <= x"0302df08";
		wait for Clk_period;
		Addr <=  "0010010000100";
		Trees_din <= x"05ff5304";
		wait for Clk_period;
		Addr <=  "0010010000101";
		Trees_din <= x"000a1245";
		wait for Clk_period;
		Addr <=  "0010010000110";
		Trees_din <= x"ffa31245";
		wait for Clk_period;
		Addr <=  "0010010000111";
		Trees_din <= x"08004104";
		wait for Clk_period;
		Addr <=  "0010010001000";
		Trees_din <= x"00b61245";
		wait for Clk_period;
		Addr <=  "0010010001001";
		Trees_din <= x"00161245";
		wait for Clk_period;
		Addr <=  "0010010001010";
		Trees_din <= x"0005f204";
		wait for Clk_period;
		Addr <=  "0010010001011";
		Trees_din <= x"ff7b1245";
		wait for Clk_period;
		Addr <=  "0010010001100";
		Trees_din <= x"ffef1245";
		wait for Clk_period;
		Addr <=  "0010010001101";
		Trees_din <= x"06d10d04";
		wait for Clk_period;
		Addr <=  "0010010001110";
		Trees_din <= x"fff31245";
		wait for Clk_period;
		Addr <=  "0010010001111";
		Trees_din <= x"00871245";
		wait for Clk_period;
		Addr <=  "0010010010000";
		Trees_din <= x"ff7a1245";
		wait for Clk_period;
		Addr <=  "0010010010001";
		Trees_din <= x"00fe360c";
		wait for Clk_period;
		Addr <=  "0010010010010";
		Trees_din <= x"18004408";
		wait for Clk_period;
		Addr <=  "0010010010011";
		Trees_din <= x"07008104";
		wait for Clk_period;
		Addr <=  "0010010010100";
		Trees_din <= x"ffaf12d1";
		wait for Clk_period;
		Addr <=  "0010010010101";
		Trees_din <= x"004f12d1";
		wait for Clk_period;
		Addr <=  "0010010010110";
		Trees_din <= x"ff6e12d1";
		wait for Clk_period;
		Addr <=  "0010010010111";
		Trees_din <= x"060aff38";
		wait for Clk_period;
		Addr <=  "0010010011000";
		Trees_din <= x"00036a1c";
		wait for Clk_period;
		Addr <=  "0010010011001";
		Trees_din <= x"1701d80c";
		wait for Clk_period;
		Addr <=  "0010010011010";
		Trees_din <= x"0b004b04";
		wait for Clk_period;
		Addr <=  "0010010011011";
		Trees_din <= x"004912d1";
		wait for Clk_period;
		Addr <=  "0010010011100";
		Trees_din <= x"00014e04";
		wait for Clk_period;
		Addr <=  "0010010011101";
		Trees_din <= x"ff6e12d1";
		wait for Clk_period;
		Addr <=  "0010010011110";
		Trees_din <= x"ffd312d1";
		wait for Clk_period;
		Addr <=  "0010010011111";
		Trees_din <= x"10023d08";
		wait for Clk_period;
		Addr <=  "0010010100000";
		Trees_din <= x"1300bd04";
		wait for Clk_period;
		Addr <=  "0010010100001";
		Trees_din <= x"000d12d1";
		wait for Clk_period;
		Addr <=  "0010010100010";
		Trees_din <= x"ffb612d1";
		wait for Clk_period;
		Addr <=  "0010010100011";
		Trees_din <= x"0a014704";
		wait for Clk_period;
		Addr <=  "0010010100100";
		Trees_din <= x"ffe212d1";
		wait for Clk_period;
		Addr <=  "0010010100101";
		Trees_din <= x"00c612d1";
		wait for Clk_period;
		Addr <=  "0010010100110";
		Trees_din <= x"08004f10";
		wait for Clk_period;
		Addr <=  "0010010100111";
		Trees_din <= x"0500a708";
		wait for Clk_period;
		Addr <=  "0010010101000";
		Trees_din <= x"07072704";
		wait for Clk_period;
		Addr <=  "0010010101001";
		Trees_din <= x"007a12d1";
		wait for Clk_period;
		Addr <=  "0010010101010";
		Trees_din <= x"002512d1";
		wait for Clk_period;
		Addr <=  "0010010101011";
		Trees_din <= x"00103e04";
		wait for Clk_period;
		Addr <=  "0010010101100";
		Trees_din <= x"ffd012d1";
		wait for Clk_period;
		Addr <=  "0010010101101";
		Trees_din <= x"005d12d1";
		wait for Clk_period;
		Addr <=  "0010010101110";
		Trees_din <= x"00079208";
		wait for Clk_period;
		Addr <=  "0010010101111";
		Trees_din <= x"05fd3604";
		wait for Clk_period;
		Addr <=  "0010010110000";
		Trees_din <= x"fff012d1";
		wait for Clk_period;
		Addr <=  "0010010110001";
		Trees_din <= x"ff8512d1";
		wait for Clk_period;
		Addr <=  "0010010110010";
		Trees_din <= x"004a12d1";
		wait for Clk_period;
		Addr <=  "0010010110011";
		Trees_din <= x"ff7d12d1";
		wait for Clk_period;
		Addr <=  "0010010110100";
		Trees_din <= x"00fe360c";
		wait for Clk_period;
		Addr <=  "0010010110101";
		Trees_din <= x"18004408";
		wait for Clk_period;
		Addr <=  "0010010110110";
		Trees_din <= x"0c012004";
		wait for Clk_period;
		Addr <=  "0010010110111";
		Trees_din <= x"fff013cd";
		wait for Clk_period;
		Addr <=  "0010010111000";
		Trees_din <= x"001913cd";
		wait for Clk_period;
		Addr <=  "0010010111001";
		Trees_din <= x"ff7013cd";
		wait for Clk_period;
		Addr <=  "0010010111010";
		Trees_din <= x"00001f34";
		wait for Clk_period;
		Addr <=  "0010010111011";
		Trees_din <= x"0a00d31c";
		wait for Clk_period;
		Addr <=  "0010010111100";
		Trees_din <= x"1604000c";
		wait for Clk_period;
		Addr <=  "0010010111101";
		Trees_din <= x"08005a08";
		wait for Clk_period;
		Addr <=  "0010010111110";
		Trees_din <= x"11000004";
		wait for Clk_period;
		Addr <=  "0010010111111";
		Trees_din <= x"005813cd";
		wait for Clk_period;
		Addr <=  "0010011000000";
		Trees_din <= x"ff8d13cd";
		wait for Clk_period;
		Addr <=  "0010011000001";
		Trees_din <= x"008a13cd";
		wait for Clk_period;
		Addr <=  "0010011000010";
		Trees_din <= x"11000008";
		wait for Clk_period;
		Addr <=  "0010011000011";
		Trees_din <= x"01fe5a04";
		wait for Clk_period;
		Addr <=  "0010011000100";
		Trees_din <= x"ff8213cd";
		wait for Clk_period;
		Addr <=  "0010011000101";
		Trees_din <= x"000413cd";
		wait for Clk_period;
		Addr <=  "0010011000110";
		Trees_din <= x"01fd3b04";
		wait for Clk_period;
		Addr <=  "0010011000111";
		Trees_din <= x"00ed13cd";
		wait for Clk_period;
		Addr <=  "0010011001000";
		Trees_din <= x"ffd413cd";
		wait for Clk_period;
		Addr <=  "0010011001001";
		Trees_din <= x"1703ac10";
		wait for Clk_period;
		Addr <=  "0010011001010";
		Trees_din <= x"0403c008";
		wait for Clk_period;
		Addr <=  "0010011001011";
		Trees_din <= x"0b00b704";
		wait for Clk_period;
		Addr <=  "0010011001100";
		Trees_din <= x"ffbc13cd";
		wait for Clk_period;
		Addr <=  "0010011001101";
		Trees_din <= x"009c13cd";
		wait for Clk_period;
		Addr <=  "0010011001110";
		Trees_din <= x"09004f04";
		wait for Clk_period;
		Addr <=  "0010011001111";
		Trees_din <= x"ffab13cd";
		wait for Clk_period;
		Addr <=  "0010011010000";
		Trees_din <= x"008413cd";
		wait for Clk_period;
		Addr <=  "0010011010001";
		Trees_din <= x"0f007a04";
		wait for Clk_period;
		Addr <=  "0010011010010";
		Trees_din <= x"002213cd";
		wait for Clk_period;
		Addr <=  "0010011010011";
		Trees_din <= x"015613cd";
		wait for Clk_period;
		Addr <=  "0010011010100";
		Trees_din <= x"12004220";
		wait for Clk_period;
		Addr <=  "0010011010101";
		Trees_din <= x"18005d10";
		wait for Clk_period;
		Addr <=  "0010011010110";
		Trees_din <= x"02fc7308";
		wait for Clk_period;
		Addr <=  "0010011010111";
		Trees_din <= x"0001c404";
		wait for Clk_period;
		Addr <=  "0010011011000";
		Trees_din <= x"ff9613cd";
		wait for Clk_period;
		Addr <=  "0010011011001";
		Trees_din <= x"001913cd";
		wait for Clk_period;
		Addr <=  "0010011011010";
		Trees_din <= x"0b00d704";
		wait for Clk_period;
		Addr <=  "0010011011011";
		Trees_din <= x"fffd13cd";
		wait for Clk_period;
		Addr <=  "0010011011100";
		Trees_din <= x"008a13cd";
		wait for Clk_period;
		Addr <=  "0010011011101";
		Trees_din <= x"10015108";
		wait for Clk_period;
		Addr <=  "0010011011110";
		Trees_din <= x"0600b904";
		wait for Clk_period;
		Addr <=  "0010011011111";
		Trees_din <= x"004713cd";
		wait for Clk_period;
		Addr <=  "0010011100000";
		Trees_din <= x"010113cd";
		wait for Clk_period;
		Addr <=  "0010011100001";
		Trees_din <= x"1702f604";
		wait for Clk_period;
		Addr <=  "0010011100010";
		Trees_din <= x"001b13cd";
		wait for Clk_period;
		Addr <=  "0010011100011";
		Trees_din <= x"000713cd";
		wait for Clk_period;
		Addr <=  "0010011100100";
		Trees_din <= x"1300ad10";
		wait for Clk_period;
		Addr <=  "0010011100101";
		Trees_din <= x"07005708";
		wait for Clk_period;
		Addr <=  "0010011100110";
		Trees_din <= x"0401c404";
		wait for Clk_period;
		Addr <=  "0010011100111";
		Trees_din <= x"ffeb13cd";
		wait for Clk_period;
		Addr <=  "0010011101000";
		Trees_din <= x"00b213cd";
		wait for Clk_period;
		Addr <=  "0010011101001";
		Trees_din <= x"1300a404";
		wait for Clk_period;
		Addr <=  "0010011101010";
		Trees_din <= x"ffde13cd";
		wait for Clk_period;
		Addr <=  "0010011101011";
		Trees_din <= x"005113cd";
		wait for Clk_period;
		Addr <=  "0010011101100";
		Trees_din <= x"02fa1a08";
		wait for Clk_period;
		Addr <=  "0010011101101";
		Trees_din <= x"01fdfe04";
		wait for Clk_period;
		Addr <=  "0010011101110";
		Trees_din <= x"ffb213cd";
		wait for Clk_period;
		Addr <=  "0010011101111";
		Trees_din <= x"00a213cd";
		wait for Clk_period;
		Addr <=  "0010011110000";
		Trees_din <= x"1e028704";
		wait for Clk_period;
		Addr <=  "0010011110001";
		Trees_din <= x"ff7e13cd";
		wait for Clk_period;
		Addr <=  "0010011110010";
		Trees_din <= x"002813cd";
		wait for Clk_period;
		Addr <=  "0010011110011";
		Trees_din <= x"00fec41c";
		wait for Clk_period;
		Addr <=  "0010011110100";
		Trees_din <= x"07008e08";
		wait for Clk_period;
		Addr <=  "0010011110101";
		Trees_din <= x"02f9d904";
		wait for Clk_period;
		Addr <=  "0010011110110";
		Trees_din <= x"000d1479";
		wait for Clk_period;
		Addr <=  "0010011110111";
		Trees_din <= x"ff6f1479";
		wait for Clk_period;
		Addr <=  "0010011111000";
		Trees_din <= x"02fb0808";
		wait for Clk_period;
		Addr <=  "0010011111001";
		Trees_din <= x"03fece04";
		wait for Clk_period;
		Addr <=  "0010011111010";
		Trees_din <= x"ff7d1479";
		wait for Clk_period;
		Addr <=  "0010011111011";
		Trees_din <= x"002d1479";
		wait for Clk_period;
		Addr <=  "0010011111100";
		Trees_din <= x"02fbc108";
		wait for Clk_period;
		Addr <=  "0010011111101";
		Trees_din <= x"11003d04";
		wait for Clk_period;
		Addr <=  "0010011111110";
		Trees_din <= x"00081479";
		wait for Clk_period;
		Addr <=  "0010011111111";
		Trees_din <= x"00b01479";
		wait for Clk_period;
		Addr <=  "0010100000000";
		Trees_din <= x"ff9f1479";
		wait for Clk_period;
		Addr <=  "0010100000001";
		Trees_din <= x"0009bd38";
		wait for Clk_period;
		Addr <=  "0010100000010";
		Trees_din <= x"01fea31c";
		wait for Clk_period;
		Addr <=  "0010100000011";
		Trees_din <= x"05ff5310";
		wait for Clk_period;
		Addr <=  "0010100000100";
		Trees_din <= x"0d006508";
		wait for Clk_period;
		Addr <=  "0010100000101";
		Trees_din <= x"16031204";
		wait for Clk_period;
		Addr <=  "0010100000110";
		Trees_din <= x"004a1479";
		wait for Clk_period;
		Addr <=  "0010100000111";
		Trees_din <= x"ffa81479";
		wait for Clk_period;
		Addr <=  "0010100001000";
		Trees_din <= x"0c027504";
		wait for Clk_period;
		Addr <=  "0010100001001";
		Trees_din <= x"002b1479";
		wait for Clk_period;
		Addr <=  "0010100001010";
		Trees_din <= x"ffb11479";
		wait for Clk_period;
		Addr <=  "0010100001011";
		Trees_din <= x"12004408";
		wait for Clk_period;
		Addr <=  "0010100001100";
		Trees_din <= x"00019e04";
		wait for Clk_period;
		Addr <=  "0010100001101";
		Trees_din <= x"ffa61479";
		wait for Clk_period;
		Addr <=  "0010100001110";
		Trees_din <= x"00381479";
		wait for Clk_period;
		Addr <=  "0010100001111";
		Trees_din <= x"ff771479";
		wait for Clk_period;
		Addr <=  "0010100010000";
		Trees_din <= x"0d00640c";
		wait for Clk_period;
		Addr <=  "0010100010001";
		Trees_din <= x"06fbc904";
		wait for Clk_period;
		Addr <=  "0010100010010";
		Trees_din <= x"ffaa1479";
		wait for Clk_period;
		Addr <=  "0010100010011";
		Trees_din <= x"09004004";
		wait for Clk_period;
		Addr <=  "0010100010100";
		Trees_din <= x"ffe81479";
		wait for Clk_period;
		Addr <=  "0010100010101";
		Trees_din <= x"00d11479";
		wait for Clk_period;
		Addr <=  "0010100010110";
		Trees_din <= x"02fda008";
		wait for Clk_period;
		Addr <=  "0010100010111";
		Trees_din <= x"070a2304";
		wait for Clk_period;
		Addr <=  "0010100011000";
		Trees_din <= x"ff691479";
		wait for Clk_period;
		Addr <=  "0010100011001";
		Trees_din <= x"000e1479";
		wait for Clk_period;
		Addr <=  "0010100011010";
		Trees_din <= x"0c01b304";
		wait for Clk_period;
		Addr <=  "0010100011011";
		Trees_din <= x"ffa11479";
		wait for Clk_period;
		Addr <=  "0010100011100";
		Trees_din <= x"00561479";
		wait for Clk_period;
		Addr <=  "0010100011101";
		Trees_din <= x"006d1479";
		wait for Clk_period;
		Addr <=  "0010100011110";
		Trees_din <= x"00fe360c";
		wait for Clk_period;
		Addr <=  "0010100011111";
		Trees_din <= x"18004408";
		wait for Clk_period;
		Addr <=  "0010100100000";
		Trees_din <= x"1f027204";
		wait for Clk_period;
		Addr <=  "0010100100001";
		Trees_din <= x"fff61505";
		wait for Clk_period;
		Addr <=  "0010100100010";
		Trees_din <= x"00121505";
		wait for Clk_period;
		Addr <=  "0010100100011";
		Trees_din <= x"ff731505";
		wait for Clk_period;
		Addr <=  "0010100100100";
		Trees_din <= x"060aff38";
		wait for Clk_period;
		Addr <=  "0010100100101";
		Trees_din <= x"0e001f18";
		wait for Clk_period;
		Addr <=  "0010100100110";
		Trees_din <= x"0e00190c";
		wait for Clk_period;
		Addr <=  "0010100100111";
		Trees_din <= x"03fe1d08";
		wait for Clk_period;
		Addr <=  "0010100101000";
		Trees_din <= x"04056704";
		wait for Clk_period;
		Addr <=  "0010100101001";
		Trees_din <= x"00781505";
		wait for Clk_period;
		Addr <=  "0010100101010";
		Trees_din <= x"ffad1505";
		wait for Clk_period;
		Addr <=  "0010100101011";
		Trees_din <= x"ffaf1505";
		wait for Clk_period;
		Addr <=  "0010100101100";
		Trees_din <= x"0002ac04";
		wait for Clk_period;
		Addr <=  "0010100101101";
		Trees_din <= x"ff6f1505";
		wait for Clk_period;
		Addr <=  "0010100101110";
		Trees_din <= x"1703d504";
		wait for Clk_period;
		Addr <=  "0010100101111";
		Trees_din <= x"ffc71505";
		wait for Clk_period;
		Addr <=  "0010100110000";
		Trees_din <= x"00251505";
		wait for Clk_period;
		Addr <=  "0010100110001";
		Trees_din <= x"09003410";
		wait for Clk_period;
		Addr <=  "0010100110010";
		Trees_din <= x"0d007708";
		wait for Clk_period;
		Addr <=  "0010100110011";
		Trees_din <= x"06034f04";
		wait for Clk_period;
		Addr <=  "0010100110100";
		Trees_din <= x"00211505";
		wait for Clk_period;
		Addr <=  "0010100110101";
		Trees_din <= x"ff9b1505";
		wait for Clk_period;
		Addr <=  "0010100110110";
		Trees_din <= x"0703b104";
		wait for Clk_period;
		Addr <=  "0010100110111";
		Trees_din <= x"00c01505";
		wait for Clk_period;
		Addr <=  "0010100111000";
		Trees_din <= x"ffe81505";
		wait for Clk_period;
		Addr <=  "0010100111001";
		Trees_din <= x"0a000408";
		wait for Clk_period;
		Addr <=  "0010100111010";
		Trees_din <= x"0403df04";
		wait for Clk_period;
		Addr <=  "0010100111011";
		Trees_din <= x"00051505";
		wait for Clk_period;
		Addr <=  "0010100111100";
		Trees_din <= x"ff6e1505";
		wait for Clk_period;
		Addr <=  "0010100111101";
		Trees_din <= x"16040004";
		wait for Clk_period;
		Addr <=  "0010100111110";
		Trees_din <= x"00031505";
		wait for Clk_period;
		Addr <=  "0010100111111";
		Trees_din <= x"00651505";
		wait for Clk_period;
		Addr <=  "0010101000000";
		Trees_din <= x"ff831505";
		wait for Clk_period;
		Addr <=  "0010101000001";
		Trees_din <= x"00fe360c";
		wait for Clk_period;
		Addr <=  "0010101000010";
		Trees_din <= x"18004408";
		wait for Clk_period;
		Addr <=  "0010101000011";
		Trees_din <= x"1703bb04";
		wait for Clk_period;
		Addr <=  "0010101000100";
		Trees_din <= x"001115b1";
		wait for Clk_period;
		Addr <=  "0010101000101";
		Trees_din <= x"fff815b1";
		wait for Clk_period;
		Addr <=  "0010101000110";
		Trees_din <= x"ff7515b1";
		wait for Clk_period;
		Addr <=  "0010101000111";
		Trees_din <= x"0003f528";
		wait for Clk_period;
		Addr <=  "0010101001000";
		Trees_din <= x"04009710";
		wait for Clk_period;
		Addr <=  "0010101001001";
		Trees_din <= x"0a02560c";
		wait for Clk_period;
		Addr <=  "0010101001010";
		Trees_din <= x"02000504";
		wait for Clk_period;
		Addr <=  "0010101001011";
		Trees_din <= x"ff6d15b1";
		wait for Clk_period;
		Addr <=  "0010101001100";
		Trees_din <= x"0303b804";
		wait for Clk_period;
		Addr <=  "0010101001101";
		Trees_din <= x"002815b1";
		wait for Clk_period;
		Addr <=  "0010101001110";
		Trees_din <= x"ff9a15b1";
		wait for Clk_period;
		Addr <=  "0010101001111";
		Trees_din <= x"004015b1";
		wait for Clk_period;
		Addr <=  "0010101010000";
		Trees_din <= x"05fb6508";
		wait for Clk_period;
		Addr <=  "0010101010001";
		Trees_din <= x"02fcf504";
		wait for Clk_period;
		Addr <=  "0010101010010";
		Trees_din <= x"ff7f15b1";
		wait for Clk_period;
		Addr <=  "0010101010011";
		Trees_din <= x"ffec15b1";
		wait for Clk_period;
		Addr <=  "0010101010100";
		Trees_din <= x"17020008";
		wait for Clk_period;
		Addr <=  "0010101010101";
		Trees_din <= x"16018204";
		wait for Clk_period;
		Addr <=  "0010101010110";
		Trees_din <= x"003b15b1";
		wait for Clk_period;
		Addr <=  "0010101010111";
		Trees_din <= x"ff7d15b1";
		wait for Clk_period;
		Addr <=  "0010101011000";
		Trees_din <= x"0a00b704";
		wait for Clk_period;
		Addr <=  "0010101011001";
		Trees_din <= x"fffb15b1";
		wait for Clk_period;
		Addr <=  "0010101011010";
		Trees_din <= x"003d15b1";
		wait for Clk_period;
		Addr <=  "0010101011011";
		Trees_din <= x"19000618";
		wait for Clk_period;
		Addr <=  "0010101011100";
		Trees_din <= x"05034010";
		wait for Clk_period;
		Addr <=  "0010101011101";
		Trees_din <= x"1300a208";
		wait for Clk_period;
		Addr <=  "0010101011110";
		Trees_din <= x"14004304";
		wait for Clk_period;
		Addr <=  "0010101011111";
		Trees_din <= x"ffdb15b1";
		wait for Clk_period;
		Addr <=  "0010101100000";
		Trees_din <= x"006715b1";
		wait for Clk_period;
		Addr <=  "0010101100001";
		Trees_din <= x"01ffbf04";
		wait for Clk_period;
		Addr <=  "0010101100010";
		Trees_din <= x"008f15b1";
		wait for Clk_period;
		Addr <=  "0010101100011";
		Trees_din <= x"001a15b1";
		wait for Clk_period;
		Addr <=  "0010101100100";
		Trees_din <= x"0c018904";
		wait for Clk_period;
		Addr <=  "0010101100101";
		Trees_din <= x"ffd015b1";
		wait for Clk_period;
		Addr <=  "0010101100110";
		Trees_din <= x"002615b1";
		wait for Clk_period;
		Addr <=  "0010101100111";
		Trees_din <= x"00079208";
		wait for Clk_period;
		Addr <=  "0010101101000";
		Trees_din <= x"18006a04";
		wait for Clk_period;
		Addr <=  "0010101101001";
		Trees_din <= x"001015b1";
		wait for Clk_period;
		Addr <=  "0010101101010";
		Trees_din <= x"ff8d15b1";
		wait for Clk_period;
		Addr <=  "0010101101011";
		Trees_din <= x"005015b1";
		wait for Clk_period;
		Addr <=  "0010101101100";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  5
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"01fe9524";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"1103e81c";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"1af84304";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"fff300d5";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"14005c10";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"08003208";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"05fe4a04";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"ff8800d5";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"003700d5";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"01fddd04";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"ff5400d5";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"ff6100d5";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"02fb0e04";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"003700d5";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"ff9000d5";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"04041504";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"00ca00d5";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"ff9000d5";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"0403251c";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"02fb570c";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"04009708";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"02fae504";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"ff9600d5";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"017b00d5";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"ff6400d5";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"15039b0c";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"04014a04";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"ff5200d5";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"05029304";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"ff5c00d5";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"00a600d5";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"000f00d5";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"01012c14";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"040b2b10";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"01ffb308";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"0609f204";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"ffdf00d5";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"ff5700d5";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"06fca304";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"ff6f00d5";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"00c200d5";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"ff5500d5";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"06f7dc10";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"040ab808";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"02019c04";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"012900d5";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"ff8800d5";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"02035104";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"ff6500d5";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"003700d5";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"18005604";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"ff9c00d5";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"031900d5";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"01fe9524";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"1103e81c";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"1af84304";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"fff801a1";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"14005c10";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"14001c08";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"10014204";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"ff9301a1";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"003701a1";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"01fddd04";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"ff5901a1";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"ff6901a1";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"09003e04";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"ff9601a1";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"004301a1";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"12004d04";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"00d601a1";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"ff9001a1";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"0403251c";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"02fb570c";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"04009708";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"02fae504";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"ff9f01a1";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"013901a1";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"ff6c01a1";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"1c06a90c";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"04014a04";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"ff5801a1";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"05029304";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"ff6201a1";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"009101a1";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"001b01a1";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"040b2b1c";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"01ffb30c";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"0609f208";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"11000004";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"00c801a1";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"ffd001a1";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"ff5d01a1";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"05fe6e08";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"01012c04";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"009c01a1";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"01df01a1";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"19000004";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"ff9001a1";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"009d01a1";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"09004804";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"ff5a01a1";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"03fc3904";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"ff8301a1";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"00ca01a1";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"01fe9530";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"1103e828";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"01fddd10";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"10030a04";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"ff5c028d";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"16025204";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"ff64028d";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"01fd1b04";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"00d1028d";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"ffa6028d";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"02f9d90c";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"05fd4508";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"00fd5304";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"015d028d";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"ffc6028d";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"ff69028d";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"08003204";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"003f028d";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"0c038704";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"ff69028d";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"0031028d";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"0c000304";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"ff93028d";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"00ce028d";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"04032520";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"02fc1010";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"04015d0c";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"01fed904";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"ff8a028d";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"04fe3e04";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"ff9b028d";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"0105028d";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"ff6f028d";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"1efbd304";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"003c028d";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"0a033004";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"ff5b028d";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"0f007004";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"0042028d";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"ff81028d";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"040b2b1c";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"01ffb30c";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"0609f208";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"08004f04";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"ffd5028d";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"008f028d";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"ff62028d";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"09004508";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"18006404";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"0032028d";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"00f8028d";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"00fca104";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"00a1028d";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"ff6e028d";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"09004804";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"ff5f028d";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"03fc3904";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"ff8c028d";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"00b9028d";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"01fe9530";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"1103e828";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"01fddd10";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"10030a04";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"ff5f0381";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"16025204";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"ff680381";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"08004104";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"00dd0381";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"ffa40381";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"02f9d90c";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"02f9d308";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"00fd5304";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"00520381";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"ff7d0381";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"00ba0381";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"08003204";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"003e0381";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"0c038704";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"ff6f0381";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"00340381";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"12004704";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"00d70381";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"ff950381";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"04032524";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"02fc1014";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"04015d10";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"19000108";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"12004304";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"003f0381";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"ff870381";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"00fdf404";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"01210381";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"00060381";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"ff760381";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"1efbd304";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"003f0381";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"0a033004";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"ff5f0381";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"0f007004";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"00400381";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"ff890381";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"040b2b1c";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"01ff9210";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"02fa6008";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"0d007c04";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"ffd50381";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"00e90381";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"17040004";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"ff9f0381";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"007c0381";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"02019c08";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"01015604";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"00460381";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"01320381";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"ff750381";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"09004804";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"ff640381";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"03fc3904";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"ff930381";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"00ac0381";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"01fe9538";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"1103e830";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"01fddd10";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"10030a04";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"ff620475";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"16025204";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"ff6c0475";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"06067c04";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"00cf0475";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"ffa60475";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"04053210";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"0f009a08";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"0e004c04";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"ff600475";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"ffd80475";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"0a01c904";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"ff9c0475";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"003f0475";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"0c028f08";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"07018e04";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"ff720475";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"ffc80475";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"15f7ba04";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"02060475";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"ffc20475";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"1cfa9c04";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"00d40475";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"ff960475";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"05fed928";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"06f84108";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"0c029a04";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"ff660475";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"001a0475";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"0701bc10";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"01002708";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"0c015104";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"ff9f0475";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"000f0475";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"00fcf104";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"010b0475";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"ffbc0475";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"1c027508";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"04082404";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"017a0475";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"001d0475";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"06fbc904";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"01320475";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"ffa80475";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"04071a10";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"1c06a90c";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"03fb8b04";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"00110475";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"1af8f804";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"fff30475";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"ff690475";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"00430475";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"03fe5804";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"ff770475";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"08004804";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"00070475";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"01210475";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"01fe9538";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"1103e830";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"01fddd10";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"10030a04";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"ff650551";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"16025204";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"ff710551";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"11007404";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"ffaa0551";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"00b60551";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"04053210";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"1f028708";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"0e004c04";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"ff620551";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"ffe20551";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"05ff4704";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"ffa50551";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"00450551";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"0c028f08";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"00fd6704";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"ffe70551";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"ff7d0551";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"15f7ba04";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"017f0551";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"ffcc0551";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"04033304";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"00c20551";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"ff9b0551";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"04fdfa04";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"ff640551";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"0609f21c";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"040b2b10";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"01ff1708";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"08005a04";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"ffd60551";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"011b0551";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"06f84104";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"ffd20551";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"00640551";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"09004804";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"ff6a0551";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"0101b404";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"ff9d0551";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"00ba0551";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"01ffcd0c";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"09004904";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"ff670551";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"12004d04";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"ffa40551";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"00400551";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"04055508";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"03fdf004";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"014e0551";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"00310551";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"ff850551";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"01fe9540";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"01fddd14";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"1103e810";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"10030a04";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"ff670625";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"16025204";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"ff750625";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"00fdde04";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"ffab0625";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"00b00625";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"00300625";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"02f9d910";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"05fc3804";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"00d10625";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"0c028f08";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"10000c04";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"002a0625";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"ff720625";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"00640625";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"01fdf40c";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"0700b404";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"ff700625";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"11000b04";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"ffaa0625";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"01220625";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"0c028808";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"0e004c04";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"ff6d0625";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"ffdc0625";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"18005d04";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"00dc0625";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"ff8b0625";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"04fdfa04";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"ff670625";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"01015614";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"06f84104";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"ff690625";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"0701bc08";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"15019e04";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"ffda0625";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"00be0625";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"0a016004";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"008d0625";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"ffa30625";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"0207e910";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"040d9708";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"0a002004";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"00270625";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"00e20625";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"1300a904";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"00400625";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"ff9f0625";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"ff990625";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"01fe5c20";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"1cfa9c08";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"0e003104";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"ffa106d1";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"00c106d1";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"13013614";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"00fb6004";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"001806d1";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"05fc3808";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"05fc3104";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"ff9106d1";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"00cd06d1";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"0c02a904";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"ff6b06d1";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"ff9306d1";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"002b06d1";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"04fdfa04";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"ff6906d1";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"0609f21c";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"040b2b10";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"11000008";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"05fddb04";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"00ca06d1";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"ff7d06d1";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"11013e04";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"fff706d1";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"008106d1";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"09004804";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"ff7006d1";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"0101b404";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"ffa706d1";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"009d06d1";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"01ffcd0c";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"09004904";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"ff6906d1";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"0402d004";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"004306d1";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"ffa706d1";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"04055508";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"02fae204";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"015806d1";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"002806d1";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"ff9206d1";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"01fe5c3c";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"1103e834";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"01fddd18";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"10030a10";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"08005608";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"03fabd04";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"ffa507d5";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"ff6607d5";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"0701d104";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"ff8407d5";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"004907d5";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"16025204";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"ff7d07d5";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"005507d5";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"18006310";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"14003708";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"17026a04";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"006707d5";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"ff6e07d5";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"19000004";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"018307d5";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"ffd007d5";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"06013008";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"09004604";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"ff8907d5";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"00d307d5";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"ff6607d5";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"12004704";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"00a807d5";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"ffac07d5";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"02fc3724";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"06f84104";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"ff7607d5";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"06038610";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"08004d08";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"08004204";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"009b07d5";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"ffd907d5";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"05fcaa04";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"001907d5";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"01ba07d5";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"09003808";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"0b008104";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"00d007d5";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"ff7407d5";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"1702f104";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"ffa507d5";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"004807d5";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"0401c408";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"1102ac04";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"ff6907d5";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"003907d5";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"0100e310";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"0b00e608";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"0e004704";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"ff7107d5";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"005e07d5";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"01ff5004";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"ff9107d5";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"008e07d5";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"02fd4d04";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"00ee07d5";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"0a008204";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"ff9907d5";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"006707d5";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"01fe5c48";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"0f008830";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"05fcae18";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"01fde808";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"0b00f504";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"ff6b08d5";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"002408d5";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"02fa3208";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"0a007204";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"ffa208d5";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"016608d5";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"11013e04";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"ff8408d5";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"001f08d5";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"10031c10";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"03fabd08";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"0d006504";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"004208d5";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"ff8608d5";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"01fe4604";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"ff6808d5";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"ffb008d5";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"05fd6f04";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"003c08d5";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"ff8f08d5";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"0700bc08";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"0c02bf04";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"ff6f08d5";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"002108d5";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"03fcda04";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"ff7e08d5";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"06088308";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"05fc5f04";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"00d608d5";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"ffa408d5";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"015708d5";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"04fdfa04";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"ff6e08d5";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"01ff1714";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"00ff2210";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"0e002f08";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"02fa6004";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"002f08d5";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"ff7808d5";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"1603fe04";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"008708d5";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"ffbf08d5";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"ff6908d5";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"08004110";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"19000008";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"0b00ed04";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"ffae08d5";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"006a08d5";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"0c020104";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"00ec08d5";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"001f08d5";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"11000008";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"0c008604";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"000408d5";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"012e08d5";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"0b006a04";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"007408d5";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"ffb308d5";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"01fe5c40";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"0f008828";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"05fcae14";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"01fde808";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"0b00f504";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"ff6d0a19";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"00230a19";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"01fe2508";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"02fa3204";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"01350a19";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"ffce0a19";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"ff880a19";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"10031c0c";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"0405b104";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"ff660a19";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"0405c504";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"00bb0a19";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"ff790a19";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"1e027a04";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"003e0a19";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"ff940a19";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"0700bc08";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"0c02bf04";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"ff720a19";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"00210a19";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"03fcda04";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"ff820a19";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"0c016a08";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"1afcad04";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"01650a19";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"00210a19";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"ffac0a19";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"02fc3740";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"1c025c20";
		wait for Clk_period;
		Addr <=  "0001001010111";
		Trees_din <= x"1b025810";
		wait for Clk_period;
		Addr <=  "0001001011000";
		Trees_din <= x"0d006c08";
		wait for Clk_period;
		Addr <=  "0001001011001";
		Trees_din <= x"0c000204";
		wait for Clk_period;
		Addr <=  "0001001011010";
		Trees_din <= x"000a0a19";
		wait for Clk_period;
		Addr <=  "0001001011011";
		Trees_din <= x"ff7a0a19";
		wait for Clk_period;
		Addr <=  "0001001011100";
		Trees_din <= x"10001b04";
		wait for Clk_period;
		Addr <=  "0001001011101";
		Trees_din <= x"00b30a19";
		wait for Clk_period;
		Addr <=  "0001001011110";
		Trees_din <= x"ffb10a19";
		wait for Clk_period;
		Addr <=  "0001001011111";
		Trees_din <= x"10003108";
		wait for Clk_period;
		Addr <=  "0001001100000";
		Trees_din <= x"04063804";
		wait for Clk_period;
		Addr <=  "0001001100001";
		Trees_din <= x"00960a19";
		wait for Clk_period;
		Addr <=  "0001001100010";
		Trees_din <= x"ff8d0a19";
		wait for Clk_period;
		Addr <=  "0001001100011";
		Trees_din <= x"0e003504";
		wait for Clk_period;
		Addr <=  "0001001100100";
		Trees_din <= x"00af0a19";
		wait for Clk_period;
		Addr <=  "0001001100101";
		Trees_din <= x"020f0a19";
		wait for Clk_period;
		Addr <=  "0001001100110";
		Trees_din <= x"1e028410";
		wait for Clk_period;
		Addr <=  "0001001100111";
		Trees_din <= x"00fd9808";
		wait for Clk_period;
		Addr <=  "0001001101000";
		Trees_din <= x"00fd5c04";
		wait for Clk_period;
		Addr <=  "0001001101001";
		Trees_din <= x"fff20a19";
		wait for Clk_period;
		Addr <=  "0001001101010";
		Trees_din <= x"01030a19";
		wait for Clk_period;
		Addr <=  "0001001101011";
		Trees_din <= x"16040004";
		wait for Clk_period;
		Addr <=  "0001001101100";
		Trees_din <= x"ff9e0a19";
		wait for Clk_period;
		Addr <=  "0001001101101";
		Trees_din <= x"008b0a19";
		wait for Clk_period;
		Addr <=  "0001001101110";
		Trees_din <= x"0c022c08";
		wait for Clk_period;
		Addr <=  "0001001101111";
		Trees_din <= x"10012c04";
		wait for Clk_period;
		Addr <=  "0001001110000";
		Trees_din <= x"ff8c0a19";
		wait for Clk_period;
		Addr <=  "0001001110001";
		Trees_din <= x"01300a19";
		wait for Clk_period;
		Addr <=  "0001001110010";
		Trees_din <= x"02fa3204";
		wait for Clk_period;
		Addr <=  "0001001110011";
		Trees_din <= x"00210a19";
		wait for Clk_period;
		Addr <=  "0001001110100";
		Trees_din <= x"ff730a19";
		wait for Clk_period;
		Addr <=  "0001001110101";
		Trees_din <= x"0401c408";
		wait for Clk_period;
		Addr <=  "0001001110110";
		Trees_din <= x"1102ac04";
		wait for Clk_period;
		Addr <=  "0001001110111";
		Trees_din <= x"ff6d0a19";
		wait for Clk_period;
		Addr <=  "0001001111000";
		Trees_din <= x"003a0a19";
		wait for Clk_period;
		Addr <=  "0001001111001";
		Trees_din <= x"00ff040c";
		wait for Clk_period;
		Addr <=  "0001001111010";
		Trees_din <= x"22000008";
		wait for Clk_period;
		Addr <=  "0001001111011";
		Trees_din <= x"06f9a104";
		wait for Clk_period;
		Addr <=  "0001001111100";
		Trees_din <= x"fff20a19";
		wait for Clk_period;
		Addr <=  "0001001111101";
		Trees_din <= x"ff6e0a19";
		wait for Clk_period;
		Addr <=  "0001001111110";
		Trees_din <= x"00540a19";
		wait for Clk_period;
		Addr <=  "0001001111111";
		Trees_din <= x"03feb208";
		wait for Clk_period;
		Addr <=  "0001010000000";
		Trees_din <= x"00056e04";
		wait for Clk_period;
		Addr <=  "0001010000001";
		Trees_din <= x"ff8b0a19";
		wait for Clk_period;
		Addr <=  "0001010000010";
		Trees_din <= x"00680a19";
		wait for Clk_period;
		Addr <=  "0001010000011";
		Trees_din <= x"0c014b04";
		wait for Clk_period;
		Addr <=  "0001010000100";
		Trees_din <= x"ff9b0a19";
		wait for Clk_period;
		Addr <=  "0001010000101";
		Trees_din <= x"01080a19";
		wait for Clk_period;
		Addr <=  "0001010000110";
		Trees_din <= x"01fe5c44";
		wait for Clk_period;
		Addr <=  "0001010000111";
		Trees_din <= x"01fddd20";
		wait for Clk_period;
		Addr <=  "0001010001000";
		Trees_din <= x"0b005d08";
		wait for Clk_period;
		Addr <=  "0001010001001";
		Trees_din <= x"10003a04";
		wait for Clk_period;
		Addr <=  "0001010001010";
		Trees_din <= x"00a10b0d";
		wait for Clk_period;
		Addr <=  "0001010001011";
		Trees_din <= x"ff890b0d";
		wait for Clk_period;
		Addr <=  "0001010001100";
		Trees_din <= x"10030a10";
		wait for Clk_period;
		Addr <=  "0001010001101";
		Trees_din <= x"03fabd08";
		wait for Clk_period;
		Addr <=  "0001010001110";
		Trees_din <= x"01fd9004";
		wait for Clk_period;
		Addr <=  "0001010001111";
		Trees_din <= x"ff8a0b0d";
		wait for Clk_period;
		Addr <=  "0001010010000";
		Trees_din <= x"00480b0d";
		wait for Clk_period;
		Addr <=  "0001010010001";
		Trees_din <= x"0b00f604";
		wait for Clk_period;
		Addr <=  "0001010010010";
		Trees_din <= x"ff660b0d";
		wait for Clk_period;
		Addr <=  "0001010010011";
		Trees_din <= x"ffb90b0d";
		wait for Clk_period;
		Addr <=  "0001010010100";
		Trees_din <= x"16025204";
		wait for Clk_period;
		Addr <=  "0001010010101";
		Trees_din <= x"ff8d0b0d";
		wait for Clk_period;
		Addr <=  "0001010010110";
		Trees_din <= x"005e0b0d";
		wait for Clk_period;
		Addr <=  "0001010010111";
		Trees_din <= x"18006314";
		wait for Clk_period;
		Addr <=  "0001010011000";
		Trees_din <= x"12003f08";
		wait for Clk_period;
		Addr <=  "0001010011001";
		Trees_din <= x"03024904";
		wait for Clk_period;
		Addr <=  "0001010011010";
		Trees_din <= x"ff760b0d";
		wait for Clk_period;
		Addr <=  "0001010011011";
		Trees_din <= x"00320b0d";
		wait for Clk_period;
		Addr <=  "0001010011100";
		Trees_din <= x"04053204";
		wait for Clk_period;
		Addr <=  "0001010011101";
		Trees_din <= x"ff940b0d";
		wait for Clk_period;
		Addr <=  "0001010011110";
		Trees_din <= x"03fbe404";
		wait for Clk_period;
		Addr <=  "0001010011111";
		Trees_din <= x"ffa00b0d";
		wait for Clk_period;
		Addr <=  "0001010100000";
		Trees_din <= x"01f40b0d";
		wait for Clk_period;
		Addr <=  "0001010100001";
		Trees_din <= x"05fca00c";
		wait for Clk_period;
		Addr <=  "0001010100010";
		Trees_din <= x"09004504";
		wait for Clk_period;
		Addr <=  "0001010100011";
		Trees_din <= x"ff8c0b0d";
		wait for Clk_period;
		Addr <=  "0001010100100";
		Trees_din <= x"01fe2504";
		wait for Clk_period;
		Addr <=  "0001010100101";
		Trees_din <= x"00c90b0d";
		wait for Clk_period;
		Addr <=  "0001010100110";
		Trees_din <= x"ffb10b0d";
		wait for Clk_period;
		Addr <=  "0001010100111";
		Trees_din <= x"ff6c0b0d";
		wait for Clk_period;
		Addr <=  "0001010101000";
		Trees_din <= x"04fdfa04";
		wait for Clk_period;
		Addr <=  "0001010101001";
		Trees_din <= x"ff740b0d";
		wait for Clk_period;
		Addr <=  "0001010101010";
		Trees_din <= x"01ff1714";
		wait for Clk_period;
		Addr <=  "0001010101011";
		Trees_din <= x"00ff2210";
		wait for Clk_period;
		Addr <=  "0001010101100";
		Trees_din <= x"0609dd08";
		wait for Clk_period;
		Addr <=  "0001010101101";
		Trees_din <= x"0406fe04";
		wait for Clk_period;
		Addr <=  "0001010101110";
		Trees_din <= x"004e0b0d";
		wait for Clk_period;
		Addr <=  "0001010101111";
		Trees_din <= x"ffc10b0d";
		wait for Clk_period;
		Addr <=  "0001010110000";
		Trees_din <= x"04009704";
		wait for Clk_period;
		Addr <=  "0001010110001";
		Trees_din <= x"00340b0d";
		wait for Clk_period;
		Addr <=  "0001010110010";
		Trees_din <= x"ff730b0d";
		wait for Clk_period;
		Addr <=  "0001010110011";
		Trees_din <= x"ff6d0b0d";
		wait for Clk_period;
		Addr <=  "0001010110100";
		Trees_din <= x"04057c10";
		wait for Clk_period;
		Addr <=  "0001010110101";
		Trees_din <= x"02fd4d08";
		wait for Clk_period;
		Addr <=  "0001010110110";
		Trees_din <= x"0f006a04";
		wait for Clk_period;
		Addr <=  "0001010110111";
		Trees_din <= x"ffab0b0d";
		wait for Clk_period;
		Addr <=  "0001010111000";
		Trees_din <= x"00b30b0d";
		wait for Clk_period;
		Addr <=  "0001010111001";
		Trees_din <= x"1001f304";
		wait for Clk_period;
		Addr <=  "0001010111010";
		Trees_din <= x"ffa90b0d";
		wait for Clk_period;
		Addr <=  "0001010111011";
		Trees_din <= x"00920b0d";
		wait for Clk_period;
		Addr <=  "0001010111100";
		Trees_din <= x"02fb8608";
		wait for Clk_period;
		Addr <=  "0001010111101";
		Trees_din <= x"02fb5704";
		wait for Clk_period;
		Addr <=  "0001010111110";
		Trees_din <= x"00180b0d";
		wait for Clk_period;
		Addr <=  "0001010111111";
		Trees_din <= x"00e60b0d";
		wait for Clk_period;
		Addr <=  "0001011000000";
		Trees_din <= x"01044c04";
		wait for Clk_period;
		Addr <=  "0001011000001";
		Trees_din <= x"ffae0b0d";
		wait for Clk_period;
		Addr <=  "0001011000010";
		Trees_din <= x"006f0b0d";
		wait for Clk_period;
		Addr <=  "0001011000011";
		Trees_din <= x"01fe5c48";
		wait for Clk_period;
		Addr <=  "0001011000100";
		Trees_din <= x"0f008830";
		wait for Clk_period;
		Addr <=  "0001011000101";
		Trees_din <= x"01fde818";
		wait for Clk_period;
		Addr <=  "0001011000110";
		Trees_din <= x"10031c10";
		wait for Clk_period;
		Addr <=  "0001011000111";
		Trees_din <= x"03fabd08";
		wait for Clk_period;
		Addr <=  "0001011001000";
		Trees_din <= x"0b00b304";
		wait for Clk_period;
		Addr <=  "0001011001001";
		Trees_din <= x"00460c19";
		wait for Clk_period;
		Addr <=  "0001011001010";
		Trees_din <= x"ff8f0c19";
		wait for Clk_period;
		Addr <=  "0001011001011";
		Trees_din <= x"0b00f604";
		wait for Clk_period;
		Addr <=  "0001011001100";
		Trees_din <= x"ff670c19";
		wait for Clk_period;
		Addr <=  "0001011001101";
		Trees_din <= x"ffbb0c19";
		wait for Clk_period;
		Addr <=  "0001011001110";
		Trees_din <= x"1e027a04";
		wait for Clk_period;
		Addr <=  "0001011001111";
		Trees_din <= x"003b0c19";
		wait for Clk_period;
		Addr <=  "0001011010000";
		Trees_din <= x"ff9e0c19";
		wait for Clk_period;
		Addr <=  "0001011010001";
		Trees_din <= x"05fcae0c";
		wait for Clk_period;
		Addr <=  "0001011010010";
		Trees_din <= x"0d007308";
		wait for Clk_period;
		Addr <=  "0001011010011";
		Trees_din <= x"0f006e04";
		wait for Clk_period;
		Addr <=  "0001011010100";
		Trees_din <= x"ffa00c19";
		wait for Clk_period;
		Addr <=  "0001011010101";
		Trees_din <= x"00c40c19";
		wait for Clk_period;
		Addr <=  "0001011010110";
		Trees_din <= x"ff910c19";
		wait for Clk_period;
		Addr <=  "0001011010111";
		Trees_din <= x"0a000708";
		wait for Clk_period;
		Addr <=  "0001011011000";
		Trees_din <= x"10003a04";
		wait for Clk_period;
		Addr <=  "0001011011001";
		Trees_din <= x"ff940c19";
		wait for Clk_period;
		Addr <=  "0001011011010";
		Trees_din <= x"00df0c19";
		wait for Clk_period;
		Addr <=  "0001011011011";
		Trees_din <= x"ff6d0c19";
		wait for Clk_period;
		Addr <=  "0001011011100";
		Trees_din <= x"0700bc08";
		wait for Clk_period;
		Addr <=  "0001011011101";
		Trees_din <= x"0406b404";
		wait for Clk_period;
		Addr <=  "0001011011110";
		Trees_din <= x"ff770c19";
		wait for Clk_period;
		Addr <=  "0001011011111";
		Trees_din <= x"00210c19";
		wait for Clk_period;
		Addr <=  "0001011100000";
		Trees_din <= x"03fcda04";
		wait for Clk_period;
		Addr <=  "0001011100001";
		Trees_din <= x"ff8b0c19";
		wait for Clk_period;
		Addr <=  "0001011100010";
		Trees_din <= x"03009508";
		wait for Clk_period;
		Addr <=  "0001011100011";
		Trees_din <= x"1c027604";
		wait for Clk_period;
		Addr <=  "0001011100100";
		Trees_din <= x"00a50c19";
		wait for Clk_period;
		Addr <=  "0001011100101";
		Trees_din <= x"ff9f0c19";
		wait for Clk_period;
		Addr <=  "0001011100110";
		Trees_din <= x"011b0c19";
		wait for Clk_period;
		Addr <=  "0001011100111";
		Trees_din <= x"03ffe524";
		wait for Clk_period;
		Addr <=  "0001011101000";
		Trees_din <= x"01012c14";
		wait for Clk_period;
		Addr <=  "0001011101001";
		Trees_din <= x"06f84104";
		wait for Clk_period;
		Addr <=  "0001011101010";
		Trees_din <= x"ff7b0c19";
		wait for Clk_period;
		Addr <=  "0001011101011";
		Trees_din <= x"07015b08";
		wait for Clk_period;
		Addr <=  "0001011101100";
		Trees_din <= x"11013e04";
		wait for Clk_period;
		Addr <=  "0001011101101";
		Trees_din <= x"ffde0c19";
		wait for Clk_period;
		Addr <=  "0001011101110";
		Trees_din <= x"005d0c19";
		wait for Clk_period;
		Addr <=  "0001011101111";
		Trees_din <= x"12004304";
		wait for Clk_period;
		Addr <=  "0001011110000";
		Trees_din <= x"ffdb0c19";
		wait for Clk_period;
		Addr <=  "0001011110001";
		Trees_din <= x"00850c19";
		wait for Clk_period;
		Addr <=  "0001011110010";
		Trees_din <= x"0a00a308";
		wait for Clk_period;
		Addr <=  "0001011110011";
		Trees_din <= x"13009b04";
		wait for Clk_period;
		Addr <=  "0001011110100";
		Trees_din <= x"001d0c19";
		wait for Clk_period;
		Addr <=  "0001011110101";
		Trees_din <= x"00bd0c19";
		wait for Clk_period;
		Addr <=  "0001011110110";
		Trees_din <= x"00fe6704";
		wait for Clk_period;
		Addr <=  "0001011110111";
		Trees_din <= x"00500c19";
		wait for Clk_period;
		Addr <=  "0001011111000";
		Trees_din <= x"ff990c19";
		wait for Clk_period;
		Addr <=  "0001011111001";
		Trees_din <= x"11000b04";
		wait for Clk_period;
		Addr <=  "0001011111010";
		Trees_din <= x"ff6b0c19";
		wait for Clk_period;
		Addr <=  "0001011111011";
		Trees_din <= x"0d007210";
		wait for Clk_period;
		Addr <=  "0001011111100";
		Trees_din <= x"17033808";
		wait for Clk_period;
		Addr <=  "0001011111101";
		Trees_din <= x"02069304";
		wait for Clk_period;
		Addr <=  "0001011111110";
		Trees_din <= x"ff8f0c19";
		wait for Clk_period;
		Addr <=  "0001011111111";
		Trees_din <= x"001b0c19";
		wait for Clk_period;
		Addr <=  "0001100000000";
		Trees_din <= x"02ff3904";
		wait for Clk_period;
		Addr <=  "0001100000001";
		Trees_din <= x"00b40c19";
		wait for Clk_period;
		Addr <=  "0001100000010";
		Trees_din <= x"ffa50c19";
		wait for Clk_period;
		Addr <=  "0001100000011";
		Trees_din <= x"0c001904";
		wait for Clk_period;
		Addr <=  "0001100000100";
		Trees_din <= x"00270c19";
		wait for Clk_period;
		Addr <=  "0001100000101";
		Trees_din <= x"ff6f0c19";
		wait for Clk_period;
		Addr <=  "0001100000110";
		Trees_din <= x"01fddd24";
		wait for Clk_period;
		Addr <=  "0001100000111";
		Trees_din <= x"0b005d08";
		wait for Clk_period;
		Addr <=  "0001100001000";
		Trees_din <= x"0401d204";
		wait for Clk_period;
		Addr <=  "0001100001001";
		Trees_din <= x"00990cfd";
		wait for Clk_period;
		Addr <=  "0001100001010";
		Trees_din <= x"ff910cfd";
		wait for Clk_period;
		Addr <=  "0001100001011";
		Trees_din <= x"0a02df14";
		wait for Clk_period;
		Addr <=  "0001100001100";
		Trees_din <= x"03fabd08";
		wait for Clk_period;
		Addr <=  "0001100001101";
		Trees_din <= x"01fd9004";
		wait for Clk_period;
		Addr <=  "0001100001110";
		Trees_din <= x"ff920cfd";
		wait for Clk_period;
		Addr <=  "0001100001111";
		Trees_din <= x"004b0cfd";
		wait for Clk_period;
		Addr <=  "0001100010000";
		Trees_din <= x"0b00f604";
		wait for Clk_period;
		Addr <=  "0001100010001";
		Trees_din <= x"ff680cfd";
		wait for Clk_period;
		Addr <=  "0001100010010";
		Trees_din <= x"0c00cf04";
		wait for Clk_period;
		Addr <=  "0001100010011";
		Trees_din <= x"ff8c0cfd";
		wait for Clk_period;
		Addr <=  "0001100010100";
		Trees_din <= x"00480cfd";
		wait for Clk_period;
		Addr <=  "0001100010101";
		Trees_din <= x"0a033004";
		wait for Clk_period;
		Addr <=  "0001100010110";
		Trees_din <= x"006f0cfd";
		wait for Clk_period;
		Addr <=  "0001100010111";
		Trees_din <= x"ff920cfd";
		wait for Clk_period;
		Addr <=  "0001100011000";
		Trees_din <= x"060a1738";
		wait for Clk_period;
		Addr <=  "0001100011001";
		Trees_din <= x"02fc3720";
		wait for Clk_period;
		Addr <=  "0001100011010";
		Trees_din <= x"07fe0a10";
		wait for Clk_period;
		Addr <=  "0001100011011";
		Trees_din <= x"12004108";
		wait for Clk_period;
		Addr <=  "0001100011100";
		Trees_din <= x"0e002b04";
		wait for Clk_period;
		Addr <=  "0001100011101";
		Trees_din <= x"002f0cfd";
		wait for Clk_period;
		Addr <=  "0001100011110";
		Trees_din <= x"01da0cfd";
		wait for Clk_period;
		Addr <=  "0001100011111";
		Trees_din <= x"0f007b04";
		wait for Clk_period;
		Addr <=  "0001100100000";
		Trees_din <= x"ffc80cfd";
		wait for Clk_period;
		Addr <=  "0001100100001";
		Trees_din <= x"00bc0cfd";
		wait for Clk_period;
		Addr <=  "0001100100010";
		Trees_din <= x"0b00ec08";
		wait for Clk_period;
		Addr <=  "0001100100011";
		Trees_din <= x"00fea104";
		wait for Clk_period;
		Addr <=  "0001100100100";
		Trees_din <= x"00390cfd";
		wait for Clk_period;
		Addr <=  "0001100100101";
		Trees_din <= x"ffda0cfd";
		wait for Clk_period;
		Addr <=  "0001100100110";
		Trees_din <= x"19001704";
		wait for Clk_period;
		Addr <=  "0001100100111";
		Trees_din <= x"ff700cfd";
		wait for Clk_period;
		Addr <=  "0001100101000";
		Trees_din <= x"00260cfd";
		wait for Clk_period;
		Addr <=  "0001100101001";
		Trees_din <= x"01ff1708";
		wait for Clk_period;
		Addr <=  "0001100101010";
		Trees_din <= x"0e004c04";
		wait for Clk_period;
		Addr <=  "0001100101011";
		Trees_din <= x"ff6e0cfd";
		wait for Clk_period;
		Addr <=  "0001100101100";
		Trees_din <= x"003c0cfd";
		wait for Clk_period;
		Addr <=  "0001100101101";
		Trees_din <= x"06063a08";
		wait for Clk_period;
		Addr <=  "0001100101110";
		Trees_din <= x"0a005604";
		wait for Clk_period;
		Addr <=  "0001100101111";
		Trees_din <= x"ff6c0cfd";
		wait for Clk_period;
		Addr <=  "0001100110000";
		Trees_din <= x"000e0cfd";
		wait for Clk_period;
		Addr <=  "0001100110001";
		Trees_din <= x"0a00c504";
		wait for Clk_period;
		Addr <=  "0001100110010";
		Trees_din <= x"00e00cfd";
		wait for Clk_period;
		Addr <=  "0001100110011";
		Trees_din <= x"ffa80cfd";
		wait for Clk_period;
		Addr <=  "0001100110100";
		Trees_din <= x"01ffcd0c";
		wait for Clk_period;
		Addr <=  "0001100110101";
		Trees_din <= x"09004904";
		wait for Clk_period;
		Addr <=  "0001100110110";
		Trees_din <= x"ff6d0cfd";
		wait for Clk_period;
		Addr <=  "0001100110111";
		Trees_din <= x"05feb804";
		wait for Clk_period;
		Addr <=  "0001100111000";
		Trees_din <= x"ffaf0cfd";
		wait for Clk_period;
		Addr <=  "0001100111001";
		Trees_din <= x"00410cfd";
		wait for Clk_period;
		Addr <=  "0001100111010";
		Trees_din <= x"04055508";
		wait for Clk_period;
		Addr <=  "0001100111011";
		Trees_din <= x"02fae204";
		wait for Clk_period;
		Addr <=  "0001100111100";
		Trees_din <= x"00e50cfd";
		wait for Clk_period;
		Addr <=  "0001100111101";
		Trees_din <= x"001b0cfd";
		wait for Clk_period;
		Addr <=  "0001100111110";
		Trees_din <= x"ffa50cfd";
		wait for Clk_period;
		Addr <=  "0001100111111";
		Trees_din <= x"01fddd24";
		wait for Clk_period;
		Addr <=  "0001101000000";
		Trees_din <= x"0b005d08";
		wait for Clk_period;
		Addr <=  "0001101000001";
		Trees_din <= x"0401d204";
		wait for Clk_period;
		Addr <=  "0001101000010";
		Trees_din <= x"008a0dd1";
		wait for Clk_period;
		Addr <=  "0001101000011";
		Trees_din <= x"ff950dd1";
		wait for Clk_period;
		Addr <=  "0001101000100";
		Trees_din <= x"0a02df14";
		wait for Clk_period;
		Addr <=  "0001101000101";
		Trees_din <= x"03fabd08";
		wait for Clk_period;
		Addr <=  "0001101000110";
		Trees_din <= x"19000204";
		wait for Clk_period;
		Addr <=  "0001101000111";
		Trees_din <= x"ff950dd1";
		wait for Clk_period;
		Addr <=  "0001101001000";
		Trees_din <= x"00490dd1";
		wait for Clk_period;
		Addr <=  "0001101001001";
		Trees_din <= x"0b00f604";
		wait for Clk_period;
		Addr <=  "0001101001010";
		Trees_din <= x"ff690dd1";
		wait for Clk_period;
		Addr <=  "0001101001011";
		Trees_din <= x"00ff6c04";
		wait for Clk_period;
		Addr <=  "0001101001100";
		Trees_din <= x"ff900dd1";
		wait for Clk_period;
		Addr <=  "0001101001101";
		Trees_din <= x"00460dd1";
		wait for Clk_period;
		Addr <=  "0001101001110";
		Trees_din <= x"0a033004";
		wait for Clk_period;
		Addr <=  "0001101001111";
		Trees_din <= x"00630dd1";
		wait for Clk_period;
		Addr <=  "0001101010000";
		Trees_din <= x"ff960dd1";
		wait for Clk_period;
		Addr <=  "0001101010001";
		Trees_din <= x"060a1730";
		wait for Clk_period;
		Addr <=  "0001101010010";
		Trees_din <= x"0d008e1c";
		wait for Clk_period;
		Addr <=  "0001101010011";
		Trees_din <= x"1300cf10";
		wait for Clk_period;
		Addr <=  "0001101010100";
		Trees_din <= x"08003d08";
		wait for Clk_period;
		Addr <=  "0001101010101";
		Trees_din <= x"02f9d904";
		wait for Clk_period;
		Addr <=  "0001101010110";
		Trees_din <= x"00440dd1";
		wait for Clk_period;
		Addr <=  "0001101010111";
		Trees_din <= x"ff770dd1";
		wait for Clk_period;
		Addr <=  "0001101011000";
		Trees_din <= x"08003f04";
		wait for Clk_period;
		Addr <=  "0001101011001";
		Trees_din <= x"00a20dd1";
		wait for Clk_period;
		Addr <=  "0001101011010";
		Trees_din <= x"00000dd1";
		wait for Clk_period;
		Addr <=  "0001101011011";
		Trees_din <= x"0f008204";
		wait for Clk_period;
		Addr <=  "0001101011100";
		Trees_din <= x"ff8d0dd1";
		wait for Clk_period;
		Addr <=  "0001101011101";
		Trees_din <= x"04071a04";
		wait for Clk_period;
		Addr <=  "0001101011110";
		Trees_din <= x"01020dd1";
		wait for Clk_period;
		Addr <=  "0001101011111";
		Trees_din <= x"ffbb0dd1";
		wait for Clk_period;
		Addr <=  "0001101100000";
		Trees_din <= x"14001c04";
		wait for Clk_period;
		Addr <=  "0001101100001";
		Trees_din <= x"006d0dd1";
		wait for Clk_period;
		Addr <=  "0001101100010";
		Trees_din <= x"08005608";
		wait for Clk_period;
		Addr <=  "0001101100011";
		Trees_din <= x"02fed304";
		wait for Clk_period;
		Addr <=  "0001101100100";
		Trees_din <= x"ff6b0dd1";
		wait for Clk_period;
		Addr <=  "0001101100101";
		Trees_din <= x"ffe60dd1";
		wait for Clk_period;
		Addr <=  "0001101100110";
		Trees_din <= x"03fcc704";
		wait for Clk_period;
		Addr <=  "0001101100111";
		Trees_din <= x"005d0dd1";
		wait for Clk_period;
		Addr <=  "0001101101000";
		Trees_din <= x"ffa40dd1";
		wait for Clk_period;
		Addr <=  "0001101101001";
		Trees_din <= x"01ffcd0c";
		wait for Clk_period;
		Addr <=  "0001101101010";
		Trees_din <= x"09004904";
		wait for Clk_period;
		Addr <=  "0001101101011";
		Trees_din <= x"ff6f0dd1";
		wait for Clk_period;
		Addr <=  "0001101101100";
		Trees_din <= x"02fb4e04";
		wait for Clk_period;
		Addr <=  "0001101101101";
		Trees_din <= x"00420dd1";
		wait for Clk_period;
		Addr <=  "0001101101110";
		Trees_din <= x"ffb10dd1";
		wait for Clk_period;
		Addr <=  "0001101101111";
		Trees_din <= x"04055508";
		wait for Clk_period;
		Addr <=  "0001101110000";
		Trees_din <= x"02fae204";
		wait for Clk_period;
		Addr <=  "0001101110001";
		Trees_din <= x"00c60dd1";
		wait for Clk_period;
		Addr <=  "0001101110010";
		Trees_din <= x"001c0dd1";
		wait for Clk_period;
		Addr <=  "0001101110011";
		Trees_din <= x"ffa90dd1";
		wait for Clk_period;
		Addr <=  "0001101110100";
		Trees_din <= x"01fddd24";
		wait for Clk_period;
		Addr <=  "0001101110101";
		Trees_din <= x"0b005d08";
		wait for Clk_period;
		Addr <=  "0001101110110";
		Trees_din <= x"10003a04";
		wait for Clk_period;
		Addr <=  "0001101110111";
		Trees_din <= x"00860ed5";
		wait for Clk_period;
		Addr <=  "0001101111000";
		Trees_din <= x"ff980ed5";
		wait for Clk_period;
		Addr <=  "0001101111001";
		Trees_din <= x"10030a14";
		wait for Clk_period;
		Addr <=  "0001101111010";
		Trees_din <= x"01fdc20c";
		wait for Clk_period;
		Addr <=  "0001101111011";
		Trees_din <= x"0b00f604";
		wait for Clk_period;
		Addr <=  "0001101111100";
		Trees_din <= x"ff6a0ed5";
		wait for Clk_period;
		Addr <=  "0001101111101";
		Trees_din <= x"03fc8b04";
		wait for Clk_period;
		Addr <=  "0001101111110";
		Trees_din <= x"004b0ed5";
		wait for Clk_period;
		Addr <=  "0001101111111";
		Trees_din <= x"ff950ed5";
		wait for Clk_period;
		Addr <=  "0001110000000";
		Trees_din <= x"00fdf604";
		wait for Clk_period;
		Addr <=  "0001110000001";
		Trees_din <= x"004c0ed5";
		wait for Clk_period;
		Addr <=  "0001110000010";
		Trees_din <= x"ff980ed5";
		wait for Clk_period;
		Addr <=  "0001110000011";
		Trees_din <= x"16025204";
		wait for Clk_period;
		Addr <=  "0001110000100";
		Trees_din <= x"ff9c0ed5";
		wait for Clk_period;
		Addr <=  "0001110000101";
		Trees_din <= x"00590ed5";
		wait for Clk_period;
		Addr <=  "0001110000110";
		Trees_din <= x"02fc3740";
		wait for Clk_period;
		Addr <=  "0001110000111";
		Trees_din <= x"06038620";
		wait for Clk_period;
		Addr <=  "0001110001000";
		Trees_din <= x"07032210";
		wait for Clk_period;
		Addr <=  "0001110001001";
		Trees_din <= x"02fb7108";
		wait for Clk_period;
		Addr <=  "0001110001010";
		Trees_din <= x"040b2b04";
		wait for Clk_period;
		Addr <=  "0001110001011";
		Trees_din <= x"00c30ed5";
		wait for Clk_period;
		Addr <=  "0001110001100";
		Trees_din <= x"ffac0ed5";
		wait for Clk_period;
		Addr <=  "0001110001101";
		Trees_din <= x"0e003304";
		wait for Clk_period;
		Addr <=  "0001110001110";
		Trees_din <= x"ff900ed5";
		wait for Clk_period;
		Addr <=  "0001110001111";
		Trees_din <= x"00270ed5";
		wait for Clk_period;
		Addr <=  "0001110010000";
		Trees_din <= x"01ff1708";
		wait for Clk_period;
		Addr <=  "0001110010001";
		Trees_din <= x"0c029a04";
		wait for Clk_period;
		Addr <=  "0001110010010";
		Trees_din <= x"ff7e0ed5";
		wait for Clk_period;
		Addr <=  "0001110010011";
		Trees_din <= x"00330ed5";
		wait for Clk_period;
		Addr <=  "0001110010100";
		Trees_din <= x"01ffa604";
		wait for Clk_period;
		Addr <=  "0001110010101";
		Trees_din <= x"00810ed5";
		wait for Clk_period;
		Addr <=  "0001110010110";
		Trees_din <= x"ffc70ed5";
		wait for Clk_period;
		Addr <=  "0001110010111";
		Trees_din <= x"0406d410";
		wait for Clk_period;
		Addr <=  "0001110011000";
		Trees_din <= x"09003808";
		wait for Clk_period;
		Addr <=  "0001110011001";
		Trees_din <= x"02fbbb04";
		wait for Clk_period;
		Addr <=  "0001110011010";
		Trees_din <= x"ff730ed5";
		wait for Clk_period;
		Addr <=  "0001110011011";
		Trees_din <= x"00590ed5";
		wait for Clk_period;
		Addr <=  "0001110011100";
		Trees_din <= x"09003e04";
		wait for Clk_period;
		Addr <=  "0001110011101";
		Trees_din <= x"009c0ed5";
		wait for Clk_period;
		Addr <=  "0001110011110";
		Trees_din <= x"fffc0ed5";
		wait for Clk_period;
		Addr <=  "0001110011111";
		Trees_din <= x"01ff2a08";
		wait for Clk_period;
		Addr <=  "0001110100000";
		Trees_din <= x"05fc3804";
		wait for Clk_period;
		Addr <=  "0001110100001";
		Trees_din <= x"00010ed5";
		wait for Clk_period;
		Addr <=  "0001110100010";
		Trees_din <= x"ff690ed5";
		wait for Clk_period;
		Addr <=  "0001110100011";
		Trees_din <= x"0a000f04";
		wait for Clk_period;
		Addr <=  "0001110100100";
		Trees_din <= x"ff930ed5";
		wait for Clk_period;
		Addr <=  "0001110100101";
		Trees_din <= x"00650ed5";
		wait for Clk_period;
		Addr <=  "0001110100110";
		Trees_din <= x"01ff1708";
		wait for Clk_period;
		Addr <=  "0001110100111";
		Trees_din <= x"0e004c04";
		wait for Clk_period;
		Addr <=  "0001110101000";
		Trees_din <= x"ff6e0ed5";
		wait for Clk_period;
		Addr <=  "0001110101001";
		Trees_din <= x"00320ed5";
		wait for Clk_period;
		Addr <=  "0001110101010";
		Trees_din <= x"04034c08";
		wait for Clk_period;
		Addr <=  "0001110101011";
		Trees_din <= x"10024d04";
		wait for Clk_period;
		Addr <=  "0001110101100";
		Trees_din <= x"ff760ed5";
		wait for Clk_period;
		Addr <=  "0001110101101";
		Trees_din <= x"003d0ed5";
		wait for Clk_period;
		Addr <=  "0001110101110";
		Trees_din <= x"0405d808";
		wait for Clk_period;
		Addr <=  "0001110101111";
		Trees_din <= x"07ff2a04";
		wait for Clk_period;
		Addr <=  "0001110110000";
		Trees_din <= x"00200ed5";
		wait for Clk_period;
		Addr <=  "0001110110001";
		Trees_din <= x"00d90ed5";
		wait for Clk_period;
		Addr <=  "0001110110010";
		Trees_din <= x"01020b04";
		wait for Clk_period;
		Addr <=  "0001110110011";
		Trees_din <= x"ff8e0ed5";
		wait for Clk_period;
		Addr <=  "0001110110100";
		Trees_din <= x"00400ed5";
		wait for Clk_period;
		Addr <=  "0001110110101";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0001110110110";
		Trees_din <= x"01fddd24";
		wait for Clk_period;
		Addr <=  "0001110110111";
		Trees_din <= x"0b005d08";
		wait for Clk_period;
		Addr <=  "0001110111000";
		Trees_din <= x"0401d204";
		wait for Clk_period;
		Addr <=  "0001110111001";
		Trees_din <= x"007b0fcd";
		wait for Clk_period;
		Addr <=  "0001110111010";
		Trees_din <= x"ff9c0fcd";
		wait for Clk_period;
		Addr <=  "0001110111011";
		Trees_din <= x"0a02df14";
		wait for Clk_period;
		Addr <=  "0001110111100";
		Trees_din <= x"03fabd08";
		wait for Clk_period;
		Addr <=  "0001110111101";
		Trees_din <= x"14004304";
		wait for Clk_period;
		Addr <=  "0001110111110";
		Trees_din <= x"ff9f0fcd";
		wait for Clk_period;
		Addr <=  "0001110111111";
		Trees_din <= x"004b0fcd";
		wait for Clk_period;
		Addr <=  "0001111000000";
		Trees_din <= x"0b00f604";
		wait for Clk_period;
		Addr <=  "0001111000001";
		Trees_din <= x"ff6b0fcd";
		wait for Clk_period;
		Addr <=  "0001111000010";
		Trees_din <= x"0a001604";
		wait for Clk_period;
		Addr <=  "0001111000011";
		Trees_din <= x"ff950fcd";
		wait for Clk_period;
		Addr <=  "0001111000100";
		Trees_din <= x"004a0fcd";
		wait for Clk_period;
		Addr <=  "0001111000101";
		Trees_din <= x"11007104";
		wait for Clk_period;
		Addr <=  "0001111000110";
		Trees_din <= x"ff9d0fcd";
		wait for Clk_period;
		Addr <=  "0001111000111";
		Trees_din <= x"00610fcd";
		wait for Clk_period;
		Addr <=  "0001111001000";
		Trees_din <= x"03ffe534";
		wait for Clk_period;
		Addr <=  "0001111001001";
		Trees_din <= x"01fecd18";
		wait for Clk_period;
		Addr <=  "0001111001010";
		Trees_din <= x"08004008";
		wait for Clk_period;
		Addr <=  "0001111001011";
		Trees_din <= x"0c02ae04";
		wait for Clk_period;
		Addr <=  "0001111001100";
		Trees_din <= x"ff710fcd";
		wait for Clk_period;
		Addr <=  "0001111001101";
		Trees_din <= x"00030fcd";
		wait for Clk_period;
		Addr <=  "0001111001110";
		Trees_din <= x"0405b108";
		wait for Clk_period;
		Addr <=  "0001111001111";
		Trees_din <= x"1b025a04";
		wait for Clk_period;
		Addr <=  "0001111010000";
		Trees_din <= x"00200fcd";
		wait for Clk_period;
		Addr <=  "0001111010001";
		Trees_din <= x"ff710fcd";
		wait for Clk_period;
		Addr <=  "0001111010010";
		Trees_din <= x"1c027e04";
		wait for Clk_period;
		Addr <=  "0001111010011";
		Trees_din <= x"006b0fcd";
		wait for Clk_period;
		Addr <=  "0001111010100";
		Trees_din <= x"ff7c0fcd";
		wait for Clk_period;
		Addr <=  "0001111010101";
		Trees_din <= x"0405170c";
		wait for Clk_period;
		Addr <=  "0001111010110";
		Trees_din <= x"1602c904";
		wait for Clk_period;
		Addr <=  "0001111010111";
		Trees_din <= x"ffac0fcd";
		wait for Clk_period;
		Addr <=  "0001111011000";
		Trees_din <= x"0d008404";
		wait for Clk_period;
		Addr <=  "0001111011001";
		Trees_din <= x"00c00fcd";
		wait for Clk_period;
		Addr <=  "0001111011010";
		Trees_din <= x"000d0fcd";
		wait for Clk_period;
		Addr <=  "0001111011011";
		Trees_din <= x"00fd9808";
		wait for Clk_period;
		Addr <=  "0001111011100";
		Trees_din <= x"1300b604";
		wait for Clk_period;
		Addr <=  "0001111011101";
		Trees_din <= x"00750fcd";
		wait for Clk_period;
		Addr <=  "0001111011110";
		Trees_din <= x"ffa80fcd";
		wait for Clk_period;
		Addr <=  "0001111011111";
		Trees_din <= x"1b028404";
		wait for Clk_period;
		Addr <=  "0001111100000";
		Trees_din <= x"ffbf0fcd";
		wait for Clk_period;
		Addr <=  "0001111100001";
		Trees_din <= x"006b0fcd";
		wait for Clk_period;
		Addr <=  "0001111100010";
		Trees_din <= x"11018218";
		wait for Clk_period;
		Addr <=  "0001111100011";
		Trees_din <= x"0f006d0c";
		wait for Clk_period;
		Addr <=  "0001111100100";
		Trees_din <= x"11000a04";
		wait for Clk_period;
		Addr <=  "0001111100101";
		Trees_din <= x"ff850fcd";
		wait for Clk_period;
		Addr <=  "0001111100110";
		Trees_din <= x"11001704";
		wait for Clk_period;
		Addr <=  "0001111100111";
		Trees_din <= x"00c10fcd";
		wait for Clk_period;
		Addr <=  "0001111101000";
		Trees_din <= x"00040fcd";
		wait for Clk_period;
		Addr <=  "0001111101001";
		Trees_din <= x"14004a08";
		wait for Clk_period;
		Addr <=  "0001111101010";
		Trees_din <= x"08003e04";
		wait for Clk_period;
		Addr <=  "0001111101011";
		Trees_din <= x"ffcf0fcd";
		wait for Clk_period;
		Addr <=  "0001111101100";
		Trees_din <= x"ff6a0fcd";
		wait for Clk_period;
		Addr <=  "0001111101101";
		Trees_din <= x"001f0fcd";
		wait for Clk_period;
		Addr <=  "0001111101110";
		Trees_din <= x"06062d04";
		wait for Clk_period;
		Addr <=  "0001111101111";
		Trees_din <= x"ffae0fcd";
		wait for Clk_period;
		Addr <=  "0001111110000";
		Trees_din <= x"1afa1804";
		wait for Clk_period;
		Addr <=  "0001111110001";
		Trees_din <= x"00c40fcd";
		wait for Clk_period;
		Addr <=  "0001111110010";
		Trees_din <= x"00150fcd";
		wait for Clk_period;
		Addr <=  "0001111110011";
		Trees_din <= x"01fdc21c";
		wait for Clk_period;
		Addr <=  "0001111110100";
		Trees_din <= x"0b005d08";
		wait for Clk_period;
		Addr <=  "0001111110101";
		Trees_din <= x"10003a04";
		wait for Clk_period;
		Addr <=  "0001111110110";
		Trees_din <= x"007f1089";
		wait for Clk_period;
		Addr <=  "0001111110111";
		Trees_din <= x"ffa41089";
		wait for Clk_period;
		Addr <=  "0001111111000";
		Trees_din <= x"10030a0c";
		wait for Clk_period;
		Addr <=  "0001111111001";
		Trees_din <= x"0b00f604";
		wait for Clk_period;
		Addr <=  "0001111111010";
		Trees_din <= x"ff6c1089";
		wait for Clk_period;
		Addr <=  "0001111111011";
		Trees_din <= x"03fc8b04";
		wait for Clk_period;
		Addr <=  "0001111111100";
		Trees_din <= x"004b1089";
		wait for Clk_period;
		Addr <=  "0001111111101";
		Trees_din <= x"ff9b1089";
		wait for Clk_period;
		Addr <=  "0001111111110";
		Trees_din <= x"00ff1d04";
		wait for Clk_period;
		Addr <=  "0001111111111";
		Trees_din <= x"ffa41089";
		wait for Clk_period;
		Addr <=  "0010000000000";
		Trees_din <= x"005a1089";
		wait for Clk_period;
		Addr <=  "0010000000001";
		Trees_din <= x"060a1734";
		wait for Clk_period;
		Addr <=  "0010000000010";
		Trees_din <= x"0d008e20";
		wait for Clk_period;
		Addr <=  "0010000000011";
		Trees_din <= x"1001d910";
		wait for Clk_period;
		Addr <=  "0010000000100";
		Trees_din <= x"05fe5d08";
		wait for Clk_period;
		Addr <=  "0010000000101";
		Trees_din <= x"0a008a04";
		wait for Clk_period;
		Addr <=  "0010000000110";
		Trees_din <= x"000d1089";
		wait for Clk_period;
		Addr <=  "0010000000111";
		Trees_din <= x"00641089";
		wait for Clk_period;
		Addr <=  "0010000001000";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "0010000001001";
		Trees_din <= x"004c1089";
		wait for Clk_period;
		Addr <=  "0010000001010";
		Trees_din <= x"ffa21089";
		wait for Clk_period;
		Addr <=  "0010000001011";
		Trees_din <= x"09004008";
		wait for Clk_period;
		Addr <=  "0010000001100";
		Trees_din <= x"03fe2504";
		wait for Clk_period;
		Addr <=  "0010000001101";
		Trees_din <= x"ffb01089";
		wait for Clk_period;
		Addr <=  "0010000001110";
		Trees_din <= x"00811089";
		wait for Clk_period;
		Addr <=  "0010000001111";
		Trees_din <= x"01020b04";
		wait for Clk_period;
		Addr <=  "0010000010000";
		Trees_din <= x"ff6c1089";
		wait for Clk_period;
		Addr <=  "0010000010001";
		Trees_din <= x"001d1089";
		wait for Clk_period;
		Addr <=  "0010000010010";
		Trees_din <= x"0a02680c";
		wait for Clk_period;
		Addr <=  "0010000010011";
		Trees_din <= x"1cfbec04";
		wait for Clk_period;
		Addr <=  "0010000010100";
		Trees_din <= x"00301089";
		wait for Clk_period;
		Addr <=  "0010000010101";
		Trees_din <= x"00009e04";
		wait for Clk_period;
		Addr <=  "0010000010110";
		Trees_din <= x"ff6f1089";
		wait for Clk_period;
		Addr <=  "0010000010111";
		Trees_din <= x"fff51089";
		wait for Clk_period;
		Addr <=  "0010000011000";
		Trees_din <= x"11000d04";
		wait for Clk_period;
		Addr <=  "0010000011001";
		Trees_din <= x"00881089";
		wait for Clk_period;
		Addr <=  "0010000011010";
		Trees_din <= x"ffe51089";
		wait for Clk_period;
		Addr <=  "0010000011011";
		Trees_din <= x"01ffcd08";
		wait for Clk_period;
		Addr <=  "0010000011100";
		Trees_din <= x"09004904";
		wait for Clk_period;
		Addr <=  "0010000011101";
		Trees_din <= x"ff721089";
		wait for Clk_period;
		Addr <=  "0010000011110";
		Trees_din <= x"fff91089";
		wait for Clk_period;
		Addr <=  "0010000011111";
		Trees_din <= x"01000904";
		wait for Clk_period;
		Addr <=  "0010000100000";
		Trees_din <= x"008c1089";
		wait for Clk_period;
		Addr <=  "0010000100001";
		Trees_din <= x"ffe91089";
		wait for Clk_period;
		Addr <=  "0010000100010";
		Trees_din <= x"01fdc218";
		wait for Clk_period;
		Addr <=  "0010000100011";
		Trees_din <= x"0700d104";
		wait for Clk_period;
		Addr <=  "0010000100100";
		Trees_din <= x"ff6f113d";
		wait for Clk_period;
		Addr <=  "0010000100101";
		Trees_din <= x"04045610";
		wait for Clk_period;
		Addr <=  "0010000100110";
		Trees_din <= x"11001404";
		wait for Clk_period;
		Addr <=  "0010000100111";
		Trees_din <= x"ff98113d";
		wait for Clk_period;
		Addr <=  "0010000101000";
		Trees_din <= x"10004704";
		wait for Clk_period;
		Addr <=  "0010000101001";
		Trees_din <= x"0130113d";
		wait for Clk_period;
		Addr <=  "0010000101010";
		Trees_din <= x"0a02df04";
		wait for Clk_period;
		Addr <=  "0010000101011";
		Trees_din <= x"ffa0113d";
		wait for Clk_period;
		Addr <=  "0010000101100";
		Trees_din <= x"007e113d";
		wait for Clk_period;
		Addr <=  "0010000101101";
		Trees_din <= x"ff78113d";
		wait for Clk_period;
		Addr <=  "0010000101110";
		Trees_din <= x"03ffe524";
		wait for Clk_period;
		Addr <=  "0010000101111";
		Trees_din <= x"02f91404";
		wait for Clk_period;
		Addr <=  "0010000110000";
		Trees_din <= x"ff7c113d";
		wait for Clk_period;
		Addr <=  "0010000110001";
		Trees_din <= x"01fecd10";
		wait for Clk_period;
		Addr <=  "0010000110010";
		Trees_din <= x"09003908";
		wait for Clk_period;
		Addr <=  "0010000110011";
		Trees_din <= x"1d01cf04";
		wait for Clk_period;
		Addr <=  "0010000110100";
		Trees_din <= x"0004113d";
		wait for Clk_period;
		Addr <=  "0010000110101";
		Trees_din <= x"ff74113d";
		wait for Clk_period;
		Addr <=  "0010000110110";
		Trees_din <= x"0a000704";
		wait for Clk_period;
		Addr <=  "0010000110111";
		Trees_din <= x"009e113d";
		wait for Clk_period;
		Addr <=  "0010000111000";
		Trees_din <= x"ffeb113d";
		wait for Clk_period;
		Addr <=  "0010000111001";
		Trees_din <= x"04051708";
		wait for Clk_period;
		Addr <=  "0010000111010";
		Trees_din <= x"16031204";
		wait for Clk_period;
		Addr <=  "0010000111011";
		Trees_din <= x"ffea113d";
		wait for Clk_period;
		Addr <=  "0010000111100";
		Trees_din <= x"0092113d";
		wait for Clk_period;
		Addr <=  "0010000111101";
		Trees_din <= x"00fd9804";
		wait for Clk_period;
		Addr <=  "0010000111110";
		Trees_din <= x"0043113d";
		wait for Clk_period;
		Addr <=  "0010000111111";
		Trees_din <= x"ffee113d";
		wait for Clk_period;
		Addr <=  "0010001000000";
		Trees_din <= x"11018218";
		wait for Clk_period;
		Addr <=  "0010001000001";
		Trees_din <= x"0f006d0c";
		wait for Clk_period;
		Addr <=  "0010001000010";
		Trees_din <= x"11000a04";
		wait for Clk_period;
		Addr <=  "0010001000011";
		Trees_din <= x"ff8c113d";
		wait for Clk_period;
		Addr <=  "0010001000100";
		Trees_din <= x"11001704";
		wait for Clk_period;
		Addr <=  "0010001000101";
		Trees_din <= x"00a3113d";
		wait for Clk_period;
		Addr <=  "0010001000110";
		Trees_din <= x"ffff113d";
		wait for Clk_period;
		Addr <=  "0010001000111";
		Trees_din <= x"14004a08";
		wait for Clk_period;
		Addr <=  "0010001001000";
		Trees_din <= x"08003e04";
		wait for Clk_period;
		Addr <=  "0010001001001";
		Trees_din <= x"ffcf113d";
		wait for Clk_period;
		Addr <=  "0010001001010";
		Trees_din <= x"ff6d113d";
		wait for Clk_period;
		Addr <=  "0010001001011";
		Trees_din <= x"001a113d";
		wait for Clk_period;
		Addr <=  "0010001001100";
		Trees_din <= x"1afa1804";
		wait for Clk_period;
		Addr <=  "0010001001101";
		Trees_din <= x"008b113d";
		wait for Clk_period;
		Addr <=  "0010001001110";
		Trees_din <= x"ffe6113d";
		wait for Clk_period;
		Addr <=  "0010001001111";
		Trees_din <= x"01fdc218";
		wait for Clk_period;
		Addr <=  "0010001010000";
		Trees_din <= x"0700d104";
		wait for Clk_period;
		Addr <=  "0010001010001";
		Trees_din <= x"ff7011d9";
		wait for Clk_period;
		Addr <=  "0010001010010";
		Trees_din <= x"04045610";
		wait for Clk_period;
		Addr <=  "0010001010011";
		Trees_din <= x"11001404";
		wait for Clk_period;
		Addr <=  "0010001010100";
		Trees_din <= x"ff9c11d9";
		wait for Clk_period;
		Addr <=  "0010001010101";
		Trees_din <= x"10004704";
		wait for Clk_period;
		Addr <=  "0010001010110";
		Trees_din <= x"010911d9";
		wait for Clk_period;
		Addr <=  "0010001010111";
		Trees_din <= x"0a02df04";
		wait for Clk_period;
		Addr <=  "0010001011000";
		Trees_din <= x"ffa411d9";
		wait for Clk_period;
		Addr <=  "0010001011001";
		Trees_din <= x"007211d9";
		wait for Clk_period;
		Addr <=  "0010001011010";
		Trees_din <= x"ff7b11d9";
		wait for Clk_period;
		Addr <=  "0010001011011";
		Trees_din <= x"060a1724";
		wait for Clk_period;
		Addr <=  "0010001011100";
		Trees_din <= x"02f91404";
		wait for Clk_period;
		Addr <=  "0010001011101";
		Trees_din <= x"ff8211d9";
		wait for Clk_period;
		Addr <=  "0010001011110";
		Trees_din <= x"02f9df10";
		wait for Clk_period;
		Addr <=  "0010001011111";
		Trees_din <= x"14003708";
		wait for Clk_period;
		Addr <=  "0010001100000";
		Trees_din <= x"19001804";
		wait for Clk_period;
		Addr <=  "0010001100001";
		Trees_din <= x"ff8711d9";
		wait for Clk_period;
		Addr <=  "0010001100010";
		Trees_din <= x"003511d9";
		wait for Clk_period;
		Addr <=  "0010001100011";
		Trees_din <= x"07ff7e04";
		wait for Clk_period;
		Addr <=  "0010001100100";
		Trees_din <= x"ffa411d9";
		wait for Clk_period;
		Addr <=  "0010001100101";
		Trees_din <= x"009a11d9";
		wait for Clk_period;
		Addr <=  "0010001100110";
		Trees_din <= x"06094f08";
		wait for Clk_period;
		Addr <=  "0010001100111";
		Trees_din <= x"01ff2204";
		wait for Clk_period;
		Addr <=  "0010001101000";
		Trees_din <= x"ffd811d9";
		wait for Clk_period;
		Addr <=  "0010001101001";
		Trees_din <= x"001611d9";
		wait for Clk_period;
		Addr <=  "0010001101010";
		Trees_din <= x"04059504";
		wait for Clk_period;
		Addr <=  "0010001101011";
		Trees_din <= x"ffc611d9";
		wait for Clk_period;
		Addr <=  "0010001101100";
		Trees_din <= x"00d711d9";
		wait for Clk_period;
		Addr <=  "0010001101101";
		Trees_din <= x"01ffcd08";
		wait for Clk_period;
		Addr <=  "0010001101110";
		Trees_din <= x"0e004204";
		wait for Clk_period;
		Addr <=  "0010001101111";
		Trees_din <= x"ff7411d9";
		wait for Clk_period;
		Addr <=  "0010001110000";
		Trees_din <= x"000011d9";
		wait for Clk_period;
		Addr <=  "0010001110001";
		Trees_din <= x"04055508";
		wait for Clk_period;
		Addr <=  "0010001110010";
		Trees_din <= x"02fae204";
		wait for Clk_period;
		Addr <=  "0010001110011";
		Trees_din <= x"009c11d9";
		wait for Clk_period;
		Addr <=  "0010001110100";
		Trees_din <= x"001611d9";
		wait for Clk_period;
		Addr <=  "0010001110101";
		Trees_din <= x"ffac11d9";
		wait for Clk_period;
		Addr <=  "0010001110110";
		Trees_din <= x"01fdc218";
		wait for Clk_period;
		Addr <=  "0010001110111";
		Trees_din <= x"00ff1808";
		wait for Clk_period;
		Addr <=  "0010001111000";
		Trees_din <= x"1affcc04";
		wait for Clk_period;
		Addr <=  "0010001111001";
		Trees_din <= x"ff711285";
		wait for Clk_period;
		Addr <=  "0010001111010";
		Trees_din <= x"fff71285";
		wait for Clk_period;
		Addr <=  "0010001111011";
		Trees_din <= x"00ff2a04";
		wait for Clk_period;
		Addr <=  "0010001111100";
		Trees_din <= x"008d1285";
		wait for Clk_period;
		Addr <=  "0010001111101";
		Trees_din <= x"05fc3808";
		wait for Clk_period;
		Addr <=  "0010001111110";
		Trees_din <= x"09003b04";
		wait for Clk_period;
		Addr <=  "0010001111111";
		Trees_din <= x"00931285";
		wait for Clk_period;
		Addr <=  "0010010000000";
		Trees_din <= x"ffad1285";
		wait for Clk_period;
		Addr <=  "0010010000001";
		Trees_din <= x"ff801285";
		wait for Clk_period;
		Addr <=  "0010010000010";
		Trees_din <= x"09004b38";
		wait for Clk_period;
		Addr <=  "0010010000011";
		Trees_din <= x"09004720";
		wait for Clk_period;
		Addr <=  "0010010000100";
		Trees_din <= x"01ff2210";
		wait for Clk_period;
		Addr <=  "0010010000101";
		Trees_din <= x"00fedc08";
		wait for Clk_period;
		Addr <=  "0010010000110";
		Trees_din <= x"0d006b04";
		wait for Clk_period;
		Addr <=  "0010010000111";
		Trees_din <= x"ff9e1285";
		wait for Clk_period;
		Addr <=  "0010010001000";
		Trees_din <= x"00191285";
		wait for Clk_period;
		Addr <=  "0010010001001";
		Trees_din <= x"04feb404";
		wait for Clk_period;
		Addr <=  "0010010001010";
		Trees_din <= x"00191285";
		wait for Clk_period;
		Addr <=  "0010010001011";
		Trees_din <= x"ff7d1285";
		wait for Clk_period;
		Addr <=  "0010010001100";
		Trees_din <= x"0d008408";
		wait for Clk_period;
		Addr <=  "0010010001101";
		Trees_din <= x"18005704";
		wait for Clk_period;
		Addr <=  "0010010001110";
		Trees_din <= x"00c21285";
		wait for Clk_period;
		Addr <=  "0010010001111";
		Trees_din <= x"00161285";
		wait for Clk_period;
		Addr <=  "0010010010000";
		Trees_din <= x"00fc3c04";
		wait for Clk_period;
		Addr <=  "0010010010001";
		Trees_din <= x"00771285";
		wait for Clk_period;
		Addr <=  "0010010010010";
		Trees_din <= x"ff9f1285";
		wait for Clk_period;
		Addr <=  "0010010010011";
		Trees_din <= x"09004808";
		wait for Clk_period;
		Addr <=  "0010010010100";
		Trees_din <= x"06fe5504";
		wait for Clk_period;
		Addr <=  "0010010010101";
		Trees_din <= x"001f1285";
		wait for Clk_period;
		Addr <=  "0010010010110";
		Trees_din <= x"011f1285";
		wait for Clk_period;
		Addr <=  "0010010010111";
		Trees_din <= x"0b006508";
		wait for Clk_period;
		Addr <=  "0010010011000";
		Trees_din <= x"0b005804";
		wait for Clk_period;
		Addr <=  "0010010011001";
		Trees_din <= x"00071285";
		wait for Clk_period;
		Addr <=  "0010010011010";
		Trees_din <= x"00c31285";
		wait for Clk_period;
		Addr <=  "0010010011011";
		Trees_din <= x"0401d204";
		wait for Clk_period;
		Addr <=  "0010010011100";
		Trees_din <= x"006f1285";
		wait for Clk_period;
		Addr <=  "0010010011101";
		Trees_din <= x"ff781285";
		wait for Clk_period;
		Addr <=  "0010010011110";
		Trees_din <= x"1300df04";
		wait for Clk_period;
		Addr <=  "0010010011111";
		Trees_din <= x"ff7e1285";
		wait for Clk_period;
		Addr <=  "0010010100000";
		Trees_din <= x"fff61285";
		wait for Clk_period;
		Addr <=  "0010010100001";
		Trees_din <= x"01fdc218";
		wait for Clk_period;
		Addr <=  "0010010100010";
		Trees_din <= x"0700d104";
		wait for Clk_period;
		Addr <=  "0010010100011";
		Trees_din <= x"ff741351";
		wait for Clk_period;
		Addr <=  "0010010100100";
		Trees_din <= x"04045610";
		wait for Clk_period;
		Addr <=  "0010010100101";
		Trees_din <= x"11001404";
		wait for Clk_period;
		Addr <=  "0010010100110";
		Trees_din <= x"ffa51351";
		wait for Clk_period;
		Addr <=  "0010010100111";
		Trees_din <= x"18006804";
		wait for Clk_period;
		Addr <=  "0010010101000";
		Trees_din <= x"ffe31351";
		wait for Clk_period;
		Addr <=  "0010010101001";
		Trees_din <= x"10004704";
		wait for Clk_period;
		Addr <=  "0010010101010";
		Trees_din <= x"01021351";
		wait for Clk_period;
		Addr <=  "0010010101011";
		Trees_din <= x"001a1351";
		wait for Clk_period;
		Addr <=  "0010010101100";
		Trees_din <= x"ff811351";
		wait for Clk_period;
		Addr <=  "0010010101101";
		Trees_din <= x"0c00e320";
		wait for Clk_period;
		Addr <=  "0010010101110";
		Trees_din <= x"1900aa1c";
		wait for Clk_period;
		Addr <=  "0010010101111";
		Trees_din <= x"01ff9210";
		wait for Clk_period;
		Addr <=  "0010010110000";
		Trees_din <= x"17040008";
		wait for Clk_period;
		Addr <=  "0010010110001";
		Trees_din <= x"03faec04";
		wait for Clk_period;
		Addr <=  "0010010110010";
		Trees_din <= x"00071351";
		wait for Clk_period;
		Addr <=  "0010010110011";
		Trees_din <= x"ff781351";
		wait for Clk_period;
		Addr <=  "0010010110100";
		Trees_din <= x"1e026504";
		wait for Clk_period;
		Addr <=  "0010010110101";
		Trees_din <= x"ff831351";
		wait for Clk_period;
		Addr <=  "0010010110110";
		Trees_din <= x"00921351";
		wait for Clk_period;
		Addr <=  "0010010110111";
		Trees_din <= x"02fd4d08";
		wait for Clk_period;
		Addr <=  "0010010111000";
		Trees_din <= x"11002304";
		wait for Clk_period;
		Addr <=  "0010010111001";
		Trees_din <= x"00571351";
		wait for Clk_period;
		Addr <=  "0010010111010";
		Trees_din <= x"ff971351";
		wait for Clk_period;
		Addr <=  "0010010111011";
		Trees_din <= x"ff8a1351";
		wait for Clk_period;
		Addr <=  "0010010111100";
		Trees_din <= x"00a61351";
		wait for Clk_period;
		Addr <=  "0010010111101";
		Trees_din <= x"1702f11c";
		wait for Clk_period;
		Addr <=  "0010010111110";
		Trees_din <= x"11001510";
		wait for Clk_period;
		Addr <=  "0010010111111";
		Trees_din <= x"05fda008";
		wait for Clk_period;
		Addr <=  "0010011000000";
		Trees_din <= x"0a02bf04";
		wait for Clk_period;
		Addr <=  "0010011000001";
		Trees_din <= x"00a71351";
		wait for Clk_period;
		Addr <=  "0010011000010";
		Trees_din <= x"ff9b1351";
		wait for Clk_period;
		Addr <=  "0010011000011";
		Trees_din <= x"0d008004";
		wait for Clk_period;
		Addr <=  "0010011000100";
		Trees_din <= x"ff871351";
		wait for Clk_period;
		Addr <=  "0010011000101";
		Trees_din <= x"00261351";
		wait for Clk_period;
		Addr <=  "0010011000110";
		Trees_din <= x"08003b04";
		wait for Clk_period;
		Addr <=  "0010011000111";
		Trees_din <= x"00921351";
		wait for Clk_period;
		Addr <=  "0010011001000";
		Trees_din <= x"09003d04";
		wait for Clk_period;
		Addr <=  "0010011001001";
		Trees_din <= x"ffe31351";
		wait for Clk_period;
		Addr <=  "0010011001010";
		Trees_din <= x"ff6d1351";
		wait for Clk_period;
		Addr <=  "0010011001011";
		Trees_din <= x"09003808";
		wait for Clk_period;
		Addr <=  "0010011001100";
		Trees_din <= x"1b024804";
		wait for Clk_period;
		Addr <=  "0010011001101";
		Trees_din <= x"001c1351";
		wait for Clk_period;
		Addr <=  "0010011001110";
		Trees_din <= x"ff771351";
		wait for Clk_period;
		Addr <=  "0010011001111";
		Trees_din <= x"12005008";
		wait for Clk_period;
		Addr <=  "0010011010000";
		Trees_din <= x"08003d04";
		wait for Clk_period;
		Addr <=  "0010011010001";
		Trees_din <= x"ffb91351";
		wait for Clk_period;
		Addr <=  "0010011010010";
		Trees_din <= x"00691351";
		wait for Clk_period;
		Addr <=  "0010011010011";
		Trees_din <= x"ff821351";
		wait for Clk_period;
		Addr <=  "0010011010100";
		Trees_din <= x"01fdc218";
		wait for Clk_period;
		Addr <=  "0010011010101";
		Trees_din <= x"00ff1808";
		wait for Clk_period;
		Addr <=  "0010011010110";
		Trees_din <= x"01fdad04";
		wait for Clk_period;
		Addr <=  "0010011010111";
		Trees_din <= x"ff74142d";
		wait for Clk_period;
		Addr <=  "0010011011000";
		Trees_din <= x"ffeb142d";
		wait for Clk_period;
		Addr <=  "0010011011001";
		Trees_din <= x"0a007d04";
		wait for Clk_period;
		Addr <=  "0010011011010";
		Trees_din <= x"ff8e142d";
		wait for Clk_period;
		Addr <=  "0010011011011";
		Trees_din <= x"09003b04";
		wait for Clk_period;
		Addr <=  "0010011011100";
		Trees_din <= x"00ab142d";
		wait for Clk_period;
		Addr <=  "0010011011101";
		Trees_din <= x"1701c004";
		wait for Clk_period;
		Addr <=  "0010011011110";
		Trees_din <= x"0019142d";
		wait for Clk_period;
		Addr <=  "0010011011111";
		Trees_din <= x"ffa2142d";
		wait for Clk_period;
		Addr <=  "0010011100000";
		Trees_din <= x"02fc3138";
		wait for Clk_period;
		Addr <=  "0010011100001";
		Trees_din <= x"00fe711c";
		wait for Clk_period;
		Addr <=  "0010011100010";
		Trees_din <= x"0a00c80c";
		wait for Clk_period;
		Addr <=  "0010011100011";
		Trees_din <= x"03f9e104";
		wait for Clk_period;
		Addr <=  "0010011100100";
		Trees_din <= x"00f1142d";
		wait for Clk_period;
		Addr <=  "0010011100101";
		Trees_din <= x"00fe5004";
		wait for Clk_period;
		Addr <=  "0010011100110";
		Trees_din <= x"ffdf142d";
		wait for Clk_period;
		Addr <=  "0010011100111";
		Trees_din <= x"0089142d";
		wait for Clk_period;
		Addr <=  "0010011101000";
		Trees_din <= x"0a01a508";
		wait for Clk_period;
		Addr <=  "0010011101001";
		Trees_din <= x"0b00e504";
		wait for Clk_period;
		Addr <=  "0010011101010";
		Trees_din <= x"00a5142d";
		wait for Clk_period;
		Addr <=  "0010011101011";
		Trees_din <= x"ffa2142d";
		wait for Clk_period;
		Addr <=  "0010011101100";
		Trees_din <= x"06049104";
		wait for Clk_period;
		Addr <=  "0010011101101";
		Trees_din <= x"0060142d";
		wait for Clk_period;
		Addr <=  "0010011101110";
		Trees_din <= x"ffc4142d";
		wait for Clk_period;
		Addr <=  "0010011101111";
		Trees_din <= x"1400380c";
		wait for Clk_period;
		Addr <=  "0010011110000";
		Trees_din <= x"18006208";
		wait for Clk_period;
		Addr <=  "0010011110001";
		Trees_din <= x"06026c04";
		wait for Clk_period;
		Addr <=  "0010011110010";
		Trees_din <= x"005c142d";
		wait for Clk_period;
		Addr <=  "0010011110011";
		Trees_din <= x"ff82142d";
		wait for Clk_period;
		Addr <=  "0010011110100";
		Trees_din <= x"00d8142d";
		wait for Clk_period;
		Addr <=  "0010011110101";
		Trees_din <= x"04040508";
		wait for Clk_period;
		Addr <=  "0010011110110";
		Trees_din <= x"0607c504";
		wait for Clk_period;
		Addr <=  "0010011110111";
		Trees_din <= x"0062142d";
		wait for Clk_period;
		Addr <=  "0010011111000";
		Trees_din <= x"ffa6142d";
		wait for Clk_period;
		Addr <=  "0010011111001";
		Trees_din <= x"06005804";
		wait for Clk_period;
		Addr <=  "0010011111010";
		Trees_din <= x"ffe7142d";
		wait for Clk_period;
		Addr <=  "0010011111011";
		Trees_din <= x"ff75142d";
		wait for Clk_period;
		Addr <=  "0010011111100";
		Trees_din <= x"01ff1708";
		wait for Clk_period;
		Addr <=  "0010011111101";
		Trees_din <= x"0e004c04";
		wait for Clk_period;
		Addr <=  "0010011111110";
		Trees_din <= x"ff76142d";
		wait for Clk_period;
		Addr <=  "0010011111111";
		Trees_din <= x"002c142d";
		wait for Clk_period;
		Addr <=  "0010100000000";
		Trees_din <= x"0a012310";
		wait for Clk_period;
		Addr <=  "0010100000001";
		Trees_din <= x"04034c08";
		wait for Clk_period;
		Addr <=  "0010100000010";
		Trees_din <= x"1e024a04";
		wait for Clk_period;
		Addr <=  "0010100000011";
		Trees_din <= x"0017142d";
		wait for Clk_period;
		Addr <=  "0010100000100";
		Trees_din <= x"ff8c142d";
		wait for Clk_period;
		Addr <=  "0010100000101";
		Trees_din <= x"0405d804";
		wait for Clk_period;
		Addr <=  "0010100000110";
		Trees_din <= x"0081142d";
		wait for Clk_period;
		Addr <=  "0010100000111";
		Trees_din <= x"fff6142d";
		wait for Clk_period;
		Addr <=  "0010100001000";
		Trees_din <= x"03045f04";
		wait for Clk_period;
		Addr <=  "0010100001001";
		Trees_din <= x"ff7e142d";
		wait for Clk_period;
		Addr <=  "0010100001010";
		Trees_din <= x"ffef142d";
		wait for Clk_period;
		Addr <=  "0010100001011";
		Trees_din <= x"01fdc218";
		wait for Clk_period;
		Addr <=  "0010100001100";
		Trees_din <= x"00ff1808";
		wait for Clk_period;
		Addr <=  "0010100001101";
		Trees_din <= x"15fd3c04";
		wait for Clk_period;
		Addr <=  "0010100001110";
		Trees_din <= x"ff7614e1";
		wait for Clk_period;
		Addr <=  "0010100001111";
		Trees_din <= x"ffef14e1";
		wait for Clk_period;
		Addr <=  "0010100010000";
		Trees_din <= x"11001404";
		wait for Clk_period;
		Addr <=  "0010100010001";
		Trees_din <= x"ff9114e1";
		wait for Clk_period;
		Addr <=  "0010100010010";
		Trees_din <= x"10004704";
		wait for Clk_period;
		Addr <=  "0010100010011";
		Trees_din <= x"00c314e1";
		wait for Clk_period;
		Addr <=  "0010100010100";
		Trees_din <= x"0a02df04";
		wait for Clk_period;
		Addr <=  "0010100010101";
		Trees_din <= x"ff9c14e1";
		wait for Clk_period;
		Addr <=  "0010100010110";
		Trees_din <= x"004714e1";
		wait for Clk_period;
		Addr <=  "0010100010111";
		Trees_din <= x"060a1734";
		wait for Clk_period;
		Addr <=  "0010100011000";
		Trees_din <= x"0d008e20";
		wait for Clk_period;
		Addr <=  "0010100011001";
		Trees_din <= x"0d006c10";
		wait for Clk_period;
		Addr <=  "0010100011010";
		Trees_din <= x"10004408";
		wait for Clk_period;
		Addr <=  "0010100011011";
		Trees_din <= x"01009f04";
		wait for Clk_period;
		Addr <=  "0010100011100";
		Trees_din <= x"ff7914e1";
		wait for Clk_period;
		Addr <=  "0010100011101";
		Trees_din <= x"003414e1";
		wait for Clk_period;
		Addr <=  "0010100011110";
		Trees_din <= x"1d027404";
		wait for Clk_period;
		Addr <=  "0010100011111";
		Trees_din <= x"004a14e1";
		wait for Clk_period;
		Addr <=  "0010100100000";
		Trees_din <= x"ffb014e1";
		wait for Clk_period;
		Addr <=  "0010100100001";
		Trees_din <= x"03004a08";
		wait for Clk_period;
		Addr <=  "0010100100010";
		Trees_din <= x"07fe5104";
		wait for Clk_period;
		Addr <=  "0010100100011";
		Trees_din <= x"008d14e1";
		wait for Clk_period;
		Addr <=  "0010100100100";
		Trees_din <= x"001e14e1";
		wait for Clk_period;
		Addr <=  "0010100100101";
		Trees_din <= x"1f027904";
		wait for Clk_period;
		Addr <=  "0010100100110";
		Trees_din <= x"ff7a14e1";
		wait for Clk_period;
		Addr <=  "0010100100111";
		Trees_din <= x"002514e1";
		wait for Clk_period;
		Addr <=  "0010100101000";
		Trees_din <= x"0a02680c";
		wait for Clk_period;
		Addr <=  "0010100101001";
		Trees_din <= x"1cfbec04";
		wait for Clk_period;
		Addr <=  "0010100101010";
		Trees_din <= x"002414e1";
		wait for Clk_period;
		Addr <=  "0010100101011";
		Trees_din <= x"09004404";
		wait for Clk_period;
		Addr <=  "0010100101100";
		Trees_din <= x"ff7914e1";
		wait for Clk_period;
		Addr <=  "0010100101101";
		Trees_din <= x"ffdf14e1";
		wait for Clk_period;
		Addr <=  "0010100101110";
		Trees_din <= x"0606de04";
		wait for Clk_period;
		Addr <=  "0010100101111";
		Trees_din <= x"ffe614e1";
		wait for Clk_period;
		Addr <=  "0010100110000";
		Trees_din <= x"006f14e1";
		wait for Clk_period;
		Addr <=  "0010100110001";
		Trees_din <= x"01ffcd08";
		wait for Clk_period;
		Addr <=  "0010100110010";
		Trees_din <= x"09004904";
		wait for Clk_period;
		Addr <=  "0010100110011";
		Trees_din <= x"ff7814e1";
		wait for Clk_period;
		Addr <=  "0010100110100";
		Trees_din <= x"000014e1";
		wait for Clk_period;
		Addr <=  "0010100110101";
		Trees_din <= x"01000904";
		wait for Clk_period;
		Addr <=  "0010100110110";
		Trees_din <= x"006814e1";
		wait for Clk_period;
		Addr <=  "0010100110111";
		Trees_din <= x"ffe614e1";
		wait for Clk_period;
		Addr <=  "0010100111000";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  6
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"020d4d30";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"02051814";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"01fae008";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"02011104";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"ff7c007d";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"00a6007d";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"02035104";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"ff51007d";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"01fe4604";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"00ca007d";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"ff65007d";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"01ff220c";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"18005104";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"00ca007d";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"13009704";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"00ca007d";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"0387007d";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"0102d20c";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"04fe6808";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"01006304";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"0037007d";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"ff8c007d";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"01f5007d";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"ff59007d";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"05157908";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"07fd2b04";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"0484007d";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"0102007d";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"06c00004";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"0037007d";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"ff62007d";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"020bd328";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"02051814";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"01fae008";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"02011104";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"ff8600e9";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"009b00e9";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"02035104";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"ff5600e9";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"0d006104";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"00bc00e9";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"ff6d00e9";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"0100630c";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"0700dd08";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"10015104";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"01b900e9";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"007d00e9";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"003000e9";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"0403ad04";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"ff6000e9";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"003800e9";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"0519b40c";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"07fec708";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"1af8f804";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"006100e9";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"01bc00e9";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"fff600e9";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"ff6700e9";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"0207e920";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"0203510c";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"01fae008";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"02011104";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"ff8e015d";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"00b2015d";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"ff5a015d";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"01ff0f0c";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"0e003608";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"12003c04";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"00a7015d";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"ff7e015d";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"0161015d";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"00fd8504";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"0039015d";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"ff65015d";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"0519b418";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"0700dd10";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"1af8f804";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"004c015d";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"0e005808";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"04050004";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"0141015d";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"0080015d";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"0078015d";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"05063404";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"003c015d";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"ff95015d";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"ff66015d";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"02051814";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"02011104";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"ff5c01c1";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"01fc5a08";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"0e003c04";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"000b01c1";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"015801c1";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"05fd8304";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"000701c1";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"ff6601c1";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"05157918";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"00103e14";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"04074e10";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"0700dd08";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"0207e904";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"007301c1";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"010001c1";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"0e002c04";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"ff8c01c1";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"009a01c1";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"ffa601c1";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"ff8001c1";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"06c00004";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"003201c1";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"ff6801c1";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"02051814";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"02011104";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"ff5e0225";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"01fc5a08";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"13009f04";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"01480225";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"00020225";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"05fd8304";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"000b0225";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"ff690225";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"0519b41c";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"00103e18";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"0700dd10";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"0207e908";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"1300a304";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"ff810225";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"00ac0225";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"0e005804";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"00da0225";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"00400225";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"18008504";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"ff830225";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"00b90225";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"ff8a0225";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"ff6d0225";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"02051814";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"02011104";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"ff600281";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"01fdaa0c";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"04ff5c04";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"ff910281";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"0e003e04";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"002f0281";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"01600281";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"ff6d0281";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"0519b418";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"000d0b14";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"04074e10";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"0700dd08";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"1af84304";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"ffde0281";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"00bc0281";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"18008504";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"ff8c0281";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"00a10281";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"ffa60281";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"ffb50281";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"ff720281";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"02051814";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"02011104";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"ff6102dd";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"01fdaa0c";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"04ff5c04";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"ff9702dd";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"08004204";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"012402dd";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"002902dd";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"ff7102dd";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"0519b418";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"0213ee10";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"0006e20c";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"1001d208";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"0306ca04";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"00a202dd";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"fffe02dd";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"ffb102dd";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"ff6302dd";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"0402a804";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"00be02dd";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"000002dd";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"ff7702dd";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"02051814";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"02011104";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"ff620339";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"01fdaa0c";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"04ff5c04";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"ff9e0339";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"0e003e04";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"00230339";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"01100339";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"ff750339";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"0519b418";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"02162714";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"0006e210";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"1001d208";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"0700dd04";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"008a0339";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"ffdb0339";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"0a005304";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"ff730339";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"00090339";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"ff6d0339";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"00b30339";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"ff7d0339";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"02011104";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"ff630391";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"0213ee20";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"0306ca10";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"0701a10c";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"04085f08";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"1001d204";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"00870391";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"ffe60391";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"ff9e0391";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"ff910391";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"01008608";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"0207e904";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"ff960391";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"00780391";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"08005104";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"ff550391";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"ffdd0391";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"0402a804";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"00a40391";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"fff60391";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"02011104";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"ff6403f5";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"0216272c";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"05053c20";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"01ff2210";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"0b00d208";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"0e004604";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"00be03f5";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"000f03f5";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"0207e904";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"ffa303f5";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"007403f5";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"12004308";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"07f9be04";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"009f03f5";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"ffff03f5";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"1300aa04";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"001403f5";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"ff4c03f5";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"18005d08";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"0306ca04";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"004603f5";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"ffb703f5";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"ff6a03f5";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"009e03f5";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"02011104";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"ff650441";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"02162720";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"05053c14";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"07f28904";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"ff8e0441";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"07fece08";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"0d00a204";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"00690441";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"ffb80441";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"05013f04";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"ff8f0441";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"00340441";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"18005d08";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"0306ca04";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"003d0441";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"ffbc0441";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"ff6e0441";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"00980441";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"02011104";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"ff6504b5";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"02162734";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"01ff801c";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"0b00d20c";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"060b1e08";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"0a000604";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"001c04b5";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"00b104b5";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"000504b5";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"05011c08";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"11000704";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"001e04b5";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"ff7604b5";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"1703b204";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"001504b5";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"006e04b5";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"0306ca10";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"0c012008";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"020bd304";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"ffe604b5";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"008804b5";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"18005f04";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"002b04b5";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"ff8704b5";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"1300bf04";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"ff6f04b5";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"fff404b5";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"009104b5";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"02011104";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"ff660511";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"02162728";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"05053c20";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"01ff8010";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"0b00d208";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"0a024e04";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"009b0511";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"ffec0511";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"05011c04";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"ffad0511";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"005c0511";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"12004308";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"07f9be04";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"008a0511";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"00040511";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"0f006f04";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"00230511";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"ff7b0511";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"19000204";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"ff760511";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"fffa0511";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"008a0511";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"02011104";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"ff660585";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"020d4d24";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"06fb660c";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"09003204";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"001f0585";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"0f006f04";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"ffed0585";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"ff720585";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"03048610";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"18006c08";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"1e027104";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"ff880585";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"005f0585";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"06096c04";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"00a90585";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"fffa0585";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"1300bb04";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"ff910585";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"002a0585";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"04e28304";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"ffc00585";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"0c024008";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"0009bd04";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"00960585";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"00160585";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"04fbca04";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"00590585";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"ffbc0585";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"02011104";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"ff6705e1";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"02162728";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"05053c20";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"04ff9e10";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"0207e908";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"001f05e1";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"ff8a05e1";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"07f73e04";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"ffcd05e1";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"008605e1";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"08004208";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"0d006b04";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"003305e1";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"00b705e1";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"0c01e204";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"ffb805e1";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"007105e1";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"18005d04";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"000205e1";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"ff7f05e1";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"008205e1";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"02011104";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"ff680655";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"02162734";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"01ff801c";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"18007310";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"0a006608";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"09003704";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"00150655";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"ff890655";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"03009504";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"fff10655";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"007c0655";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"0d006004";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"00090655";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"14004704";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"00a20655";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"002f0655";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"0c01d810";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"020bd308";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"06fb6604";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"ff890655";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"000d0655";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"0a000604";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"fff20655";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"00680655";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"19000204";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"ff770655";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"ffe90655";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"007c0655";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"02011104";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"ff6806cd";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"020bd324";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"06fb6608";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"0208f904";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"ff8806cd";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"ffe006cd";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"0b00c910";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"04fdab08";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"0c00f504";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"003b06cd";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"ffb006cd";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"08004204";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"00ae06cd";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"003a06cd";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"0f006c04";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"004a06cd";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"09003c04";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"ffe506cd";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"ff8406cd";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"0c023608";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"0009bd04";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"008906cd";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"000406cd";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"17029b04";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"004706cd";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"0f007704";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"ff9106cd";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"ffe306cd";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"02011104";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"ff690729";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"02162728";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"01ff8018";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"0b00d20c";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"060b1e08";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"01fba504";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"00010729";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"00860729";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"fffb0729";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"0207e904";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"ffb30729";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"1afc4504";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"ffe70729";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"006b0729";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"00020f0c";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"0d006d04";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"ffa90729";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"12004504";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"00540729";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"ffdb0729";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"ff9f0729";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"00730729";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"02011104";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"ff690795";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"020bd324";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"01fd5910";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"0a015b0c";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"0b00c608";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"11002e04";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"00200795";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"00920795";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"00100795";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"ffe10795";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"05fdeb08";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"1603ff04";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"ffda0795";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"00660795";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"22000e08";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"0c002104";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"ffec0795";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"ff820795";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"002a0795";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"0c023608";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"0009bd04";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"00810795";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"00000795";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"17029b04";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"00400795";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"ffae0795";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"02011104";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"ff6a07f1";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"02162728";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"01ff8014";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"06053308";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"0a000604";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"ffe607f1";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"007407f1";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"1b025504";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"005807f1";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"0e003604";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"ff9307f1";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"002707f1";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"0306ca10";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"0c00cd08";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"1afc7204";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"006007f1";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"ffec07f1";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"19000104";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"ffa807f1";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"000907f1";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"ffa107f1";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"006b07f1";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"02011104";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"ff6b084d";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"0207e914";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"04ff9e08";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"12003e04";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"fff5084d";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"ff9a084d";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"08004204";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"006c084d";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"0c01e204";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"ff9e084d";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"004d084d";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"0c024010";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"03014208";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"0b00d704";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"ffd3084d";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"0038084d";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"0309a404";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"007f084d";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"000a084d";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"1e027604";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"ffbd084d";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"0030084d";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"02011104";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"ff6c08b1";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"0213ee28";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"01ff2214";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"0e00370c";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"1afcdf08";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"06030404";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"002208b1";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"ff9a08b1";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"004c08b1";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"0e004204";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"006f08b1";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"000208b1";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"09003a08";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"08004204";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"003d08b1";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"ffe008b1";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"020bd304";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"ff9208b1";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"07f5f204";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"ffae08b1";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"002e08b1";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"11007804";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"006708b1";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"001408b1";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"02011104";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"ff6d090d";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"0207e914";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"04ff9e08";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"12003e04";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"fff5090d";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"ffa1090d";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"01fc5a04";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"0062090d";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"07fa3404";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"0045090d";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"ffa2090d";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"0c024010";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"03018608";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"0e002a04";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"ffda090d";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"0035090d";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"0309a404";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"007a090d";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"000b090d";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"1e026c04";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"ffca090d";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"000e090d";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"02011104";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"ff6e0959";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"02162720";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"01ff8014";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"06053308";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"0b00e304";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"005f0959";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"00010959";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"1b025504";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"00460959";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"0e003604";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"ffa30959";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"00170959";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"18005f04";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"00190959";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"0f006f04";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"000c0959";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"ff960959";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"005d0959";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  7
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"0702cf74";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"07009b40";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"07ff5520";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"07fdaa10";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"11033508";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"01fae004";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"ffc10185";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"ff560185";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"05fe0f04";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"00ca0185";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"ff6f0185";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"0d00b308";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"0a03b804";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"ff720185";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"00150185";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"03fe6304";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"ff810185";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"00df0185";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"02faef10";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"09004b08";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"00fc3c04";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"fff80185";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"ff5a0185";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"03fcc104";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"ff790185";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"015c0185";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"01fe8c08";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"15f76004";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"00480185";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"ffc40185";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"1c023d04";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"000f0185";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"ff580185";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"04074220";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"07018e10";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"06095d08";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"1dfdbd04";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"02350185";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"00330185";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"19000304";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"ff5a0185";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"000d0185";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"00fd3408";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"0a001204";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"ffde0185";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"02e10185";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"06075004";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"01030185";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"00450185";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"0409320c";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"10036008";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"1603eb04";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"ff5d0185";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"00180185";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"01b00185";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"02fe1804";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"ff560185";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"00210185";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"0408fa2c";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"0705d21c";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"0003ad10";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"0406be08";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"0607fe04";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"02850185";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"00390185";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"00ffa104";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"012b0185";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"fff70185";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"19000808";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"0a01ac04";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"ff6a0185";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"00370185";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"012b0185";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"0009bd08";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"1e028704";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"03c20185";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"00a60185";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"05029304";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"ff740185";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"015c0185";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"07079b1c";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"0e004010";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"0e002408";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"06fdaa04";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"ffbf0185";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"01d20185";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"0c000a04";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"00370185";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"ff660185";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"02fb1608";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"00fe0604";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"ffa40185";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"00370185";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"02350185";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"13009f04";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"00a60185";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"03050185";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"07015b60";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"07ff9134";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"07fdaa18";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"11033510";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"01fae008";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"11002e04";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"ff9302e9";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"003802e9";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"0f008204";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"ff5702e9";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"ff7902e9";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"05fe0f04";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"00bb02e9";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"ff7902e9";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"0a03b810";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"0d00b308";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"05fe5d04";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"ff7002e9";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"ff9d02e9";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"09002c04";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"ff8602e9";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"00be02e9";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"05fe3e08";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"1c027504";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"004002e9";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"ff8702e9";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"013c02e9";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"05053c1c";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"1f028810";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"03fda808";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"0c030804";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"ff9602e9";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"005102e9";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"0c00a004";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"006802e9";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"ffc302e9";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"11015708";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"08004104";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"003002e9";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"025b02e9";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"ff9c02e9";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"0c003a04";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"ff9a02e9";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"0a005804";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"027602e9";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"10012f04";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"ffa902e9";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"00d602e9";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"07049c38";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"0407ad1c";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"00fd370c";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"0c000804";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"ff9202e9";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"03006f04";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"01d702e9";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"fffc02e9";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"0003f508";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"19000604";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"00cf02e9";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"001f02e9";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"0703df04";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"ff6602e9";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"004102e9";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"040a4410";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"1d027608";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"0e002904";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"005202e9";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"ff7f02e9";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"19000004";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"017f02e9";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"fff602e9";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"14002e04";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"002f02e9";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"0e004804";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"ff5c02e9";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"002102e9";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"040e5418";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"0009bd10";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"05fbbf08";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"12004c04";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"009a02e9";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"01c102e9";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"0d006c04";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"012702e9";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"01c802e9";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"0104e104";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"ff7302e9";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"014402e9";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"ff7102e9";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"07015b60";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"07ff9134";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"07fdaa18";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"11033510";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"01fc3108";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"0e001e04";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"0079045d";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"ff7b045d";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"15f6f904";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"ffaf045d";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"ff5c045d";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"05fe0f04";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"00a6045d";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"ff80045d";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"0a03b810";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"03fc7f08";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"00ff0804";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"ff5b045d";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"ffce045d";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"08005604";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"ff96045d";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"0026045d";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"11000504";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"0105045d";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"11002104";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"ff8c045d";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"003f045d";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"05043c1c";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"1f028810";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"03fda808";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"0c030804";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"ffa2045d";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"0048045d";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"0c00a004";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"005a045d";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"ffc9045d";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"0a006604";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"ffa2045d";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"0e003204";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"01bc045d";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"0029045d";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"0b00e208";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"14004404";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"ff87045d";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"00cd045d";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"11000504";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"ffa8045d";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"01d3045d";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"0703c530";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"0407ad14";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"0003f510";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"02fc7908";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"08004504";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"0033045d";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"00a5045d";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"0b007f04";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"ffc4045d";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"0164045d";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"ff6f045d";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"1afc4510";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"13009808";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"02fb5a04";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"0007045d";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"01d0045d";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"12003f04";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"004f045d";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"ff78045d";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"12004008";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"02fa8a04";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"ff83045d";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"0041045d";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"ff61045d";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"040bfb1c";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"05fd4910";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"0705d208";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"06ffea04";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"ffdd045d";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"00c4045d";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"0005f204";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"0124045d";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"000f045d";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"08003a04";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"ff80045d";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"00103e04";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"0147045d";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"ff9e045d";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"070a230c";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"05ff2208";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"1001d904";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"ff66045d";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"0038045d";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"003d045d";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"00fd045d";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"07009b50";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"07fdaa20";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"1e024210";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"04e87804";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"00b905a9";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"11033504";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"ff6a05a9";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"05fe7404";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"00d105a9";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"ffab05a9";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"01fc310c";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"00ffbd08";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"04f7bd04";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"004105a9";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"ff6c05a9";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"008c05a9";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"ff6005a9";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"05fbe914";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"03ffdb0c";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"10005808";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"0c009604";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"ff8705a9";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"01eb05a9";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"ff6f05a9";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"01fe0104";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"01f805a9";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"002405a9";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"02fbce10";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"01fd4a08";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"0d006904";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"006205a9";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"ff8205a9";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"15f71104";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"000205a9";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"ff7105a9";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"02fbd204";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"016905a9";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"0a036704";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"ffc305a9";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"00b005a9";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"07035730";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"04093220";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"03fda810";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"1d026b08";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"0a01a504";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"ffbd05a9";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"009805a9";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"07031004";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"004205a9";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"013d05a9";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"0a01bd08";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"02f96704";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"ff6e05a9";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"00a605a9";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"12004e04";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"ff8805a9";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"008205a9";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"02fe180c";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"0a022f04";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"ff6205a9";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"09004204";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"004205a9";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"ffa805a9";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"004405a9";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"040d2320";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"07072710";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"06002808";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"13007f04";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"011705a9";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"002005a9";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"1d022a04";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"ffc105a9";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"00cf05a9";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"05fb0208";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"00036a04";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"008705a9";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"ff8305a9";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"0009bd04";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"010705a9";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"001a05a9";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"1001d904";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"ff7305a9";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"003505a9";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"07009b54";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"07fdaa20";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"1e024210";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"14003b0c";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"08004708";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"02ff3904";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"ff8906ed";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"003b06ed";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"013906ed";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"ff7106ed";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"01fc310c";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"0a019f08";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"00ffbd04";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"ff7106ed";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"003c06ed";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"008d06ed";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"ff6306ed";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"01fe9520";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"02fadc10";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"0b006f08";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"03fd9a04";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"ffaa06ed";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"00f506ed";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"05febf04";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"ff6506ed";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"ffe606ed";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"07ff5508";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"0f006e04";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"002e06ed";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"ff9b06ed";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"060a9904";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"003a06ed";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"ffb606ed";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"09004b0c";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"08003c08";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"11000704";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"00d706ed";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"ff8b06ed";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"ff6506ed";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"12004804";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"009b06ed";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"ff8f06ed";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"0703572c";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"04093220";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"0d007210";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"1f027f08";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"22000004";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"ffd906ed";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"011806ed";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"04044d04";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"011206ed";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"000c06ed";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"00fd1c08";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"02fb5704";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"005706ed";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"016506ed";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"0404a804";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"007806ed";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"001706ed";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"0a000104";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"003b06ed";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"0603f604";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"ff6606ed";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"fffe06ed";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"040e5420";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"05fe2710";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"00036a08";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"01fe7c04";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"009b06ed";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"001406ed";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"070be104";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"ffd006ed";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"00da06ed";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"1300c508";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"04036d04";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"00b406ed";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"013f06ed";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"10008804";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"ff7206ed";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"009c06ed";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"ff7d06ed";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"07009b5c";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"07fdaa28";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"1e024210";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"14003b0c";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"19001308";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"08004604";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"00190829";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"01620829";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"ff8d0829";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"ff760829";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"01fc310c";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"0e001e04";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"00960829";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"09004704";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"ff750829";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"00420829";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"00fc5608";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"0f008304";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"ff7c0829";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"00460829";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"ff620829";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"01fe951c";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"02fadc10";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"06066c08";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"09004604";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"ffb10829";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"011d0829";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"05fe9704";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"ff610829";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"fff50829";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"0a03da08";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"07ff9104";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"ffc60829";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"001f0829";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"011d0829";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"09004b10";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"08003c08";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"11000604";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"00d30829";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"ff8e0829";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"07fe2104";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"ffa60829";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"ff620829";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"0b005c04";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"ff930829";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"008e0829";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"07072724";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"040c5820";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"09003410";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"0d00ab08";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"0701a104";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"fffa0829";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"00e80829";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"14002e04";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"ff520829";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"00c80829";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"0e004508";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"12004304";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"00490829";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"00050829";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"01fe7904";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"00b00829";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"ffc30829";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"ff6c0829";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"13007508";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"0f005304";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"00700829";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"ff6b0829";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"05fb0208";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"00036a04";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"00690829";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"ff960829";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"03fb0708";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"0c020a04";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"00b50829";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"ffdd0829";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"02f88d04";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"004e0829";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"00de0829";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"07015b70";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"07ff5538";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"07fdaa18";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"1800550c";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"12003f08";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"18005404";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"ff8609bd";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"003409bd";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"010109bd";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"01fae004";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"002109bd";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"15f6f904";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"ffda09bd";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"ff6309bd";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"1e026110";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"10000008";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"08004b04";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"ffa809bd";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"00c509bd";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"0a016304";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"ff6409bd";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"ffc809bd";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"15f79c08";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"0a005c04";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"ff8609bd";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"011909bd";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"0d006704";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"004709bd";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"ffa909bd";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"1b024b18";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"03fbfe08";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"16016404";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"004009bd";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"ff7009bd";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"01fd8908";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"02fc5704";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"ffb509bd";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"010a09bd";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"0f008504";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"010a09bd";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"ff9309bd";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"21000010";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"00fcd108";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"11000304";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"013f09bd";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"fff109bd";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"03031e04";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"ffbb09bd";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"007709bd";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"0607a908";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"06053304";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"ffaa09bd";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"01df09bd";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"0e001e04";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"004309bd";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"ff9b09bd";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"07072738";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"0900341c";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"08004010";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"0f007f08";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"19003104";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"ff5809bd";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"fff109bd";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"03fbba04";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"014009bd";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"004b09bd";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"14002a04";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"ff6709bd";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"02f9c104";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"001709bd";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"00f409bd";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"040a1510";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"1702d708";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"1af9e504";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"ffc509bd";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"008109bd";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"05fe2d04";
		wait for Clk_period;
		Addr <=  "0001001010111";
		Trees_din <= x"000609bd";
		wait for Clk_period;
		Addr <=  "0001001011000";
		Trees_din <= x"006209bd";
		wait for Clk_period;
		Addr <=  "0001001011001";
		Trees_din <= x"0a000104";
		wait for Clk_period;
		Addr <=  "0001001011010";
		Trees_din <= x"00ca09bd";
		wait for Clk_period;
		Addr <=  "0001001011011";
		Trees_din <= x"0e004104";
		wait for Clk_period;
		Addr <=  "0001001011100";
		Trees_din <= x"ff6709bd";
		wait for Clk_period;
		Addr <=  "0001001011101";
		Trees_din <= x"005309bd";
		wait for Clk_period;
		Addr <=  "0001001011110";
		Trees_din <= x"13007508";
		wait for Clk_period;
		Addr <=  "0001001011111";
		Trees_din <= x"0f005304";
		wait for Clk_period;
		Addr <=  "0001001100000";
		Trees_din <= x"006409bd";
		wait for Clk_period;
		Addr <=  "0001001100001";
		Trees_din <= x"ff7409bd";
		wait for Clk_period;
		Addr <=  "0001001100010";
		Trees_din <= x"00036a0c";
		wait for Clk_period;
		Addr <=  "0001001100011";
		Trees_din <= x"02f8bf08";
		wait for Clk_period;
		Addr <=  "0001001100100";
		Trees_din <= x"07094904";
		wait for Clk_period;
		Addr <=  "0001001100101";
		Trees_din <= x"ff7e09bd";
		wait for Clk_period;
		Addr <=  "0001001100110";
		Trees_din <= x"00b709bd";
		wait for Clk_period;
		Addr <=  "0001001100111";
		Trees_din <= x"00cb09bd";
		wait for Clk_period;
		Addr <=  "0001001101000";
		Trees_din <= x"1c027d08";
		wait for Clk_period;
		Addr <=  "0001001101001";
		Trees_din <= x"08004204";
		wait for Clk_period;
		Addr <=  "0001001101010";
		Trees_din <= x"002b09bd";
		wait for Clk_period;
		Addr <=  "0001001101011";
		Trees_din <= x"00ca09bd";
		wait for Clk_period;
		Addr <=  "0001001101100";
		Trees_din <= x"070be104";
		wait for Clk_period;
		Addr <=  "0001001101101";
		Trees_din <= x"ff8a09bd";
		wait for Clk_period;
		Addr <=  "0001001101110";
		Trees_din <= x"007a09bd";
		wait for Clk_period;
		Addr <=  "0001001101111";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0001001110000";
		Trees_din <= x"07009b58";
		wait for Clk_period;
		Addr <=  "0001001110001";
		Trees_din <= x"07fdaa20";
		wait for Clk_period;
		Addr <=  "0001001110010";
		Trees_din <= x"18005510";
		wait for Clk_period;
		Addr <=  "0001001110011";
		Trees_din <= x"12003f0c";
		wait for Clk_period;
		Addr <=  "0001001110100";
		Trees_din <= x"02ff3904";
		wait for Clk_period;
		Addr <=  "0001001110101";
		Trees_din <= x"ff750b5d";
		wait for Clk_period;
		Addr <=  "0001001110110";
		Trees_din <= x"01fdd904";
		wait for Clk_period;
		Addr <=  "0001001110111";
		Trees_din <= x"00a00b5d";
		wait for Clk_period;
		Addr <=  "0001001111000";
		Trees_din <= x"ff910b5d";
		wait for Clk_period;
		Addr <=  "0001001111001";
		Trees_din <= x"00d20b5d";
		wait for Clk_period;
		Addr <=  "0001001111010";
		Trees_din <= x"15f6f908";
		wait for Clk_period;
		Addr <=  "0001001111011";
		Trees_din <= x"05157904";
		wait for Clk_period;
		Addr <=  "0001001111100";
		Trees_din <= x"ff820b5d";
		wait for Clk_period;
		Addr <=  "0001001111101";
		Trees_din <= x"00c90b5d";
		wait for Clk_period;
		Addr <=  "0001001111110";
		Trees_din <= x"01fae004";
		wait for Clk_period;
		Addr <=  "0001001111111";
		Trees_din <= x"00240b5d";
		wait for Clk_period;
		Addr <=  "0001010000000";
		Trees_din <= x"ff650b5d";
		wait for Clk_period;
		Addr <=  "0001010000001";
		Trees_din <= x"01fe9520";
		wait for Clk_period;
		Addr <=  "0001010000010";
		Trees_din <= x"02fadc10";
		wait for Clk_period;
		Addr <=  "0001010000011";
		Trees_din <= x"0b006f08";
		wait for Clk_period;
		Addr <=  "0001010000100";
		Trees_din <= x"0b006104";
		wait for Clk_period;
		Addr <=  "0001010000101";
		Trees_din <= x"ffbe0b5d";
		wait for Clk_period;
		Addr <=  "0001010000110";
		Trees_din <= x"01000b5d";
		wait for Clk_period;
		Addr <=  "0001010000111";
		Trees_din <= x"05febf04";
		wait for Clk_period;
		Addr <=  "0001010001000";
		Trees_din <= x"ff6e0b5d";
		wait for Clk_period;
		Addr <=  "0001010001001";
		Trees_din <= x"00000b5d";
		wait for Clk_period;
		Addr <=  "0001010001010";
		Trees_din <= x"0d008b08";
		wait for Clk_period;
		Addr <=  "0001010001011";
		Trees_din <= x"0d006804";
		wait for Clk_period;
		Addr <=  "0001010001100";
		Trees_din <= x"004c0b5d";
		wait for Clk_period;
		Addr <=  "0001010001101";
		Trees_din <= x"ffd00b5d";
		wait for Clk_period;
		Addr <=  "0001010001110";
		Trees_din <= x"18005e04";
		wait for Clk_period;
		Addr <=  "0001010001111";
		Trees_din <= x"00da0b5d";
		wait for Clk_period;
		Addr <=  "0001010010000";
		Trees_din <= x"ff770b5d";
		wait for Clk_period;
		Addr <=  "0001010010001";
		Trees_din <= x"09004b10";
		wait for Clk_period;
		Addr <=  "0001010010010";
		Trees_din <= x"08003c08";
		wait for Clk_period;
		Addr <=  "0001010010011";
		Trees_din <= x"11000604";
		wait for Clk_period;
		Addr <=  "0001010010100";
		Trees_din <= x"00a70b5d";
		wait for Clk_period;
		Addr <=  "0001010010101";
		Trees_din <= x"ff980b5d";
		wait for Clk_period;
		Addr <=  "0001010010110";
		Trees_din <= x"07fe2104";
		wait for Clk_period;
		Addr <=  "0001010010111";
		Trees_din <= x"ffb70b5d";
		wait for Clk_period;
		Addr <=  "0001010011000";
		Trees_din <= x"ff650b5d";
		wait for Clk_period;
		Addr <=  "0001010011001";
		Trees_din <= x"12004804";
		wait for Clk_period;
		Addr <=  "0001010011010";
		Trees_din <= x"00970b5d";
		wait for Clk_period;
		Addr <=  "0001010011011";
		Trees_din <= x"ff9d0b5d";
		wait for Clk_period;
		Addr <=  "0001010011100";
		Trees_din <= x"07047c40";
		wait for Clk_period;
		Addr <=  "0001010011101";
		Trees_din <= x"00fe7120";
		wait for Clk_period;
		Addr <=  "0001010011110";
		Trees_din <= x"12004910";
		wait for Clk_period;
		Addr <=  "0001010011111";
		Trees_din <= x"21000008";
		wait for Clk_period;
		Addr <=  "0001010100000";
		Trees_din <= x"03fe4f04";
		wait for Clk_period;
		Addr <=  "0001010100001";
		Trees_din <= x"ffe70b5d";
		wait for Clk_period;
		Addr <=  "0001010100010";
		Trees_din <= x"00590b5d";
		wait for Clk_period;
		Addr <=  "0001010100011";
		Trees_din <= x"18006204";
		wait for Clk_period;
		Addr <=  "0001010100100";
		Trees_din <= x"01440b5d";
		wait for Clk_period;
		Addr <=  "0001010100101";
		Trees_din <= x"000b0b5d";
		wait for Clk_period;
		Addr <=  "0001010100110";
		Trees_din <= x"07019808";
		wait for Clk_period;
		Addr <=  "0001010100111";
		Trees_din <= x"01fd8104";
		wait for Clk_period;
		Addr <=  "0001010101000";
		Trees_din <= x"ff8a0b5d";
		wait for Clk_period;
		Addr <=  "0001010101001";
		Trees_din <= x"00870b5d";
		wait for Clk_period;
		Addr <=  "0001010101010";
		Trees_din <= x"01fe5c04";
		wait for Clk_period;
		Addr <=  "0001010101011";
		Trees_din <= x"00e80b5d";
		wait for Clk_period;
		Addr <=  "0001010101100";
		Trees_din <= x"001b0b5d";
		wait for Clk_period;
		Addr <=  "0001010101101";
		Trees_din <= x"12004410";
		wait for Clk_period;
		Addr <=  "0001010101110";
		Trees_din <= x"20040008";
		wait for Clk_period;
		Addr <=  "0001010101111";
		Trees_din <= x"0a000b04";
		wait for Clk_period;
		Addr <=  "0001010110000";
		Trees_din <= x"00790b5d";
		wait for Clk_period;
		Addr <=  "0001010110001";
		Trees_din <= x"ff8e0b5d";
		wait for Clk_period;
		Addr <=  "0001010110010";
		Trees_din <= x"03fb1704";
		wait for Clk_period;
		Addr <=  "0001010110011";
		Trees_din <= x"ffb30b5d";
		wait for Clk_period;
		Addr <=  "0001010110100";
		Trees_din <= x"007e0b5d";
		wait for Clk_period;
		Addr <=  "0001010110101";
		Trees_din <= x"10032908";
		wait for Clk_period;
		Addr <=  "0001010110110";
		Trees_din <= x"04064c04";
		wait for Clk_period;
		Addr <=  "0001010110111";
		Trees_din <= x"ffef0b5d";
		wait for Clk_period;
		Addr <=  "0001010111000";
		Trees_din <= x"ff720b5d";
		wait for Clk_period;
		Addr <=  "0001010111001";
		Trees_din <= x"05fdf504";
		wait for Clk_period;
		Addr <=  "0001010111010";
		Trees_din <= x"00ce0b5d";
		wait for Clk_period;
		Addr <=  "0001010111011";
		Trees_din <= x"ffa10b5d";
		wait for Clk_period;
		Addr <=  "0001010111100";
		Trees_din <= x"10019220";
		wait for Clk_period;
		Addr <=  "0001010111101";
		Trees_din <= x"03fb2510";
		wait for Clk_period;
		Addr <=  "0001010111110";
		Trees_din <= x"07062508";
		wait for Clk_period;
		Addr <=  "0001010111111";
		Trees_din <= x"02fbd204";
		wait for Clk_period;
		Addr <=  "0001011000000";
		Trees_din <= x"ff3f0b5d";
		wait for Clk_period;
		Addr <=  "0001011000001";
		Trees_din <= x"00530b5d";
		wait for Clk_period;
		Addr <=  "0001011000010";
		Trees_din <= x"06fd2b04";
		wait for Clk_period;
		Addr <=  "0001011000011";
		Trees_din <= x"00160b5d";
		wait for Clk_period;
		Addr <=  "0001011000100";
		Trees_din <= x"00c50b5d";
		wait for Clk_period;
		Addr <=  "0001011000101";
		Trees_din <= x"0f008708";
		wait for Clk_period;
		Addr <=  "0001011000110";
		Trees_din <= x"08004604";
		wait for Clk_period;
		Addr <=  "0001011000111";
		Trees_din <= x"00490b5d";
		wait for Clk_period;
		Addr <=  "0001011001000";
		Trees_din <= x"00c00b5d";
		wait for Clk_period;
		Addr <=  "0001011001001";
		Trees_din <= x"01fdc804";
		wait for Clk_period;
		Addr <=  "0001011001010";
		Trees_din <= x"00700b5d";
		wait for Clk_period;
		Addr <=  "0001011001011";
		Trees_din <= x"ff870b5d";
		wait for Clk_period;
		Addr <=  "0001011001100";
		Trees_din <= x"00056e10";
		wait for Clk_period;
		Addr <=  "0001011001101";
		Trees_din <= x"09004308";
		wait for Clk_period;
		Addr <=  "0001011001110";
		Trees_din <= x"0409b104";
		wait for Clk_period;
		Addr <=  "0001011001111";
		Trees_din <= x"01040b5d";
		wait for Clk_period;
		Addr <=  "0001011010000";
		Trees_din <= x"004f0b5d";
		wait for Clk_period;
		Addr <=  "0001011010001";
		Trees_din <= x"0406cb04";
		wait for Clk_period;
		Addr <=  "0001011010010";
		Trees_din <= x"00b90b5d";
		wait for Clk_period;
		Addr <=  "0001011010011";
		Trees_din <= x"ffbf0b5d";
		wait for Clk_period;
		Addr <=  "0001011010100";
		Trees_din <= x"08004004";
		wait for Clk_period;
		Addr <=  "0001011010101";
		Trees_din <= x"006b0b5d";
		wait for Clk_period;
		Addr <=  "0001011010110";
		Trees_din <= x"ff760b5d";
		wait for Clk_period;
		Addr <=  "0001011010111";
		Trees_din <= x"07ff9848";
		wait for Clk_period;
		Addr <=  "0001011011000";
		Trees_din <= x"01fe482c";
		wait for Clk_period;
		Addr <=  "0001011011001";
		Trees_din <= x"01fe251c";
		wait for Clk_period;
		Addr <=  "0001011011010";
		Trees_din <= x"0d00ae10";
		wait for Clk_period;
		Addr <=  "0001011011011";
		Trees_din <= x"0f006e08";
		wait for Clk_period;
		Addr <=  "0001011011100";
		Trees_din <= x"0e003504";
		wait for Clk_period;
		Addr <=  "0001011011101";
		Trees_din <= x"013c0c91";
		wait for Clk_period;
		Addr <=  "0001011011110";
		Trees_din <= x"ffaa0c91";
		wait for Clk_period;
		Addr <=  "0001011011111";
		Trees_din <= x"17009f04";
		wait for Clk_period;
		Addr <=  "0001011100000";
		Trees_din <= x"007e0c91";
		wait for Clk_period;
		Addr <=  "0001011100001";
		Trees_din <= x"ff990c91";
		wait for Clk_period;
		Addr <=  "0001011100010";
		Trees_din <= x"18004104";
		wait for Clk_period;
		Addr <=  "0001011100011";
		Trees_din <= x"ffab0c91";
		wait for Clk_period;
		Addr <=  "0001011100100";
		Trees_din <= x"14002a04";
		wait for Clk_period;
		Addr <=  "0001011100101";
		Trees_din <= x"015e0c91";
		wait for Clk_period;
		Addr <=  "0001011100110";
		Trees_din <= x"00210c91";
		wait for Clk_period;
		Addr <=  "0001011100111";
		Trees_din <= x"09004408";
		wait for Clk_period;
		Addr <=  "0001011101000";
		Trees_din <= x"0e001e04";
		wait for Clk_period;
		Addr <=  "0001011101001";
		Trees_din <= x"00bf0c91";
		wait for Clk_period;
		Addr <=  "0001011101010";
		Trees_din <= x"ff830c91";
		wait for Clk_period;
		Addr <=  "0001011101011";
		Trees_din <= x"02fbe704";
		wait for Clk_period;
		Addr <=  "0001011101100";
		Trees_din <= x"ffae0c91";
		wait for Clk_period;
		Addr <=  "0001011101101";
		Trees_din <= x"02e90c91";
		wait for Clk_period;
		Addr <=  "0001011101110";
		Trees_din <= x"00fd3110";
		wait for Clk_period;
		Addr <=  "0001011101111";
		Trees_din <= x"0306ca0c";
		wait for Clk_period;
		Addr <=  "0001011110000";
		Trees_din <= x"12005708";
		wait for Clk_period;
		Addr <=  "0001011110001";
		Trees_din <= x"19000804";
		wait for Clk_period;
		Addr <=  "0001011110010";
		Trees_din <= x"ff710c91";
		wait for Clk_period;
		Addr <=  "0001011110011";
		Trees_din <= x"00010c91";
		wait for Clk_period;
		Addr <=  "0001011110100";
		Trees_din <= x"003f0c91";
		wait for Clk_period;
		Addr <=  "0001011110101";
		Trees_din <= x"00eb0c91";
		wait for Clk_period;
		Addr <=  "0001011110110";
		Trees_din <= x"11000008";
		wait for Clk_period;
		Addr <=  "0001011110111";
		Trees_din <= x"11000004";
		wait for Clk_period;
		Addr <=  "0001011111000";
		Trees_din <= x"ff790c91";
		wait for Clk_period;
		Addr <=  "0001011111001";
		Trees_din <= x"00b60c91";
		wait for Clk_period;
		Addr <=  "0001011111010";
		Trees_din <= x"ff650c91";
		wait for Clk_period;
		Addr <=  "0001011111011";
		Trees_din <= x"07037220";
		wait for Clk_period;
		Addr <=  "0001011111100";
		Trees_din <= x"02f91404";
		wait for Clk_period;
		Addr <=  "0001011111101";
		Trees_din <= x"ff520c91";
		wait for Clk_period;
		Addr <=  "0001011111110";
		Trees_din <= x"04093210";
		wait for Clk_period;
		Addr <=  "0001011111111";
		Trees_din <= x"1d026b08";
		wait for Clk_period;
		Addr <=  "0001100000000";
		Trees_din <= x"1afc5704";
		wait for Clk_period;
		Addr <=  "0001100000001";
		Trees_din <= x"ff670c91";
		wait for Clk_period;
		Addr <=  "0001100000010";
		Trees_din <= x"00100c91";
		wait for Clk_period;
		Addr <=  "0001100000011";
		Trees_din <= x"1b026f04";
		wait for Clk_period;
		Addr <=  "0001100000100";
		Trees_din <= x"00bd0c91";
		wait for Clk_period;
		Addr <=  "0001100000101";
		Trees_din <= x"00200c91";
		wait for Clk_period;
		Addr <=  "0001100000110";
		Trees_din <= x"07028104";
		wait for Clk_period;
		Addr <=  "0001100000111";
		Trees_din <= x"ff6d0c91";
		wait for Clk_period;
		Addr <=  "0001100001000";
		Trees_din <= x"0e002404";
		wait for Clk_period;
		Addr <=  "0001100001001";
		Trees_din <= x"009c0c91";
		wait for Clk_period;
		Addr <=  "0001100001010";
		Trees_din <= x"ff930c91";
		wait for Clk_period;
		Addr <=  "0001100001011";
		Trees_din <= x"10019220";
		wait for Clk_period;
		Addr <=  "0001100001100";
		Trees_din <= x"11000110";
		wait for Clk_period;
		Addr <=  "0001100001101";
		Trees_din <= x"00ffb608";
		wait for Clk_period;
		Addr <=  "0001100001110";
		Trees_din <= x"1afd9004";
		wait for Clk_period;
		Addr <=  "0001100001111";
		Trees_din <= x"00fe0c91";
		wait for Clk_period;
		Addr <=  "0001100010000";
		Trees_din <= x"00250c91";
		wait for Clk_period;
		Addr <=  "0001100010001";
		Trees_din <= x"03fb7b04";
		wait for Clk_period;
		Addr <=  "0001100010010";
		Trees_din <= x"ffe00c91";
		wait for Clk_period;
		Addr <=  "0001100010011";
		Trees_din <= x"008c0c91";
		wait for Clk_period;
		Addr <=  "0001100010100";
		Trees_din <= x"1d026708";
		wait for Clk_period;
		Addr <=  "0001100010101";
		Trees_din <= x"07079b04";
		wait for Clk_period;
		Addr <=  "0001100010110";
		Trees_din <= x"ffc40c91";
		wait for Clk_period;
		Addr <=  "0001100010111";
		Trees_din <= x"00570c91";
		wait for Clk_period;
		Addr <=  "0001100011000";
		Trees_din <= x"1afb2404";
		wait for Clk_period;
		Addr <=  "0001100011001";
		Trees_din <= x"fffd0c91";
		wait for Clk_period;
		Addr <=  "0001100011010";
		Trees_din <= x"00690c91";
		wait for Clk_period;
		Addr <=  "0001100011011";
		Trees_din <= x"0c02dd0c";
		wait for Clk_period;
		Addr <=  "0001100011100";
		Trees_din <= x"09003b04";
		wait for Clk_period;
		Addr <=  "0001100011101";
		Trees_din <= x"01020c91";
		wait for Clk_period;
		Addr <=  "0001100011110";
		Trees_din <= x"0d006504";
		wait for Clk_period;
		Addr <=  "0001100011111";
		Trees_din <= x"00e90c91";
		wait for Clk_period;
		Addr <=  "0001100100000";
		Trees_din <= x"002b0c91";
		wait for Clk_period;
		Addr <=  "0001100100001";
		Trees_din <= x"0706c604";
		wait for Clk_period;
		Addr <=  "0001100100010";
		Trees_din <= x"ff710c91";
		wait for Clk_period;
		Addr <=  "0001100100011";
		Trees_din <= x"00690c91";
		wait for Clk_period;
		Addr <=  "0001100100100";
		Trees_din <= x"07ff9148";
		wait for Clk_period;
		Addr <=  "0001100100101";
		Trees_din <= x"01fe482c";
		wait for Clk_period;
		Addr <=  "0001100100110";
		Trees_din <= x"01fe2920";
		wait for Clk_period;
		Addr <=  "0001100100111";
		Trees_din <= x"060b7710";
		wait for Clk_period;
		Addr <=  "0001100101000";
		Trees_din <= x"09003608";
		wait for Clk_period;
		Addr <=  "0001100101001";
		Trees_din <= x"09003404";
		wait for Clk_period;
		Addr <=  "0001100101010";
		Trees_din <= x"ffd80e0d";
		wait for Clk_period;
		Addr <=  "0001100101011";
		Trees_din <= x"01840e0d";
		wait for Clk_period;
		Addr <=  "0001100101100";
		Trees_din <= x"060ab304";
		wait for Clk_period;
		Addr <=  "0001100101101";
		Trees_din <= x"ffac0e0d";
		wait for Clk_period;
		Addr <=  "0001100101110";
		Trees_din <= x"005e0e0d";
		wait for Clk_period;
		Addr <=  "0001100101111";
		Trees_din <= x"14002e08";
		wait for Clk_period;
		Addr <=  "0001100110000";
		Trees_din <= x"1e027004";
		wait for Clk_period;
		Addr <=  "0001100110001";
		Trees_din <= x"00d90e0d";
		wait for Clk_period;
		Addr <=  "0001100110010";
		Trees_din <= x"ff9e0e0d";
		wait for Clk_period;
		Addr <=  "0001100110011";
		Trees_din <= x"0c02f204";
		wait for Clk_period;
		Addr <=  "0001100110100";
		Trees_din <= x"ff690e0d";
		wait for Clk_period;
		Addr <=  "0001100110101";
		Trees_din <= x"003e0e0d";
		wait for Clk_period;
		Addr <=  "0001100110110";
		Trees_din <= x"12004804";
		wait for Clk_period;
		Addr <=  "0001100110111";
		Trees_din <= x"ff8a0e0d";
		wait for Clk_period;
		Addr <=  "0001100111000";
		Trees_din <= x"14004604";
		wait for Clk_period;
		Addr <=  "0001100111001";
		Trees_din <= x"01d80e0d";
		wait for Clk_period;
		Addr <=  "0001100111010";
		Trees_din <= x"00220e0d";
		wait for Clk_period;
		Addr <=  "0001100111011";
		Trees_din <= x"00fd3110";
		wait for Clk_period;
		Addr <=  "0001100111100";
		Trees_din <= x"0306ca0c";
		wait for Clk_period;
		Addr <=  "0001100111101";
		Trees_din <= x"05fed504";
		wait for Clk_period;
		Addr <=  "0001100111110";
		Trees_din <= x"ff770e0d";
		wait for Clk_period;
		Addr <=  "0001100111111";
		Trees_din <= x"03fee504";
		wait for Clk_period;
		Addr <=  "0001101000000";
		Trees_din <= x"00c80e0d";
		wait for Clk_period;
		Addr <=  "0001101000001";
		Trees_din <= x"ff8e0e0d";
		wait for Clk_period;
		Addr <=  "0001101000010";
		Trees_din <= x"00c10e0d";
		wait for Clk_period;
		Addr <=  "0001101000011";
		Trees_din <= x"11000008";
		wait for Clk_period;
		Addr <=  "0001101000100";
		Trees_din <= x"11000004";
		wait for Clk_period;
		Addr <=  "0001101000101";
		Trees_din <= x"ff7f0e0d";
		wait for Clk_period;
		Addr <=  "0001101000110";
		Trees_din <= x"009f0e0d";
		wait for Clk_period;
		Addr <=  "0001101000111";
		Trees_din <= x"ff670e0d";
		wait for Clk_period;
		Addr <=  "0001101001000";
		Trees_din <= x"07018e3c";
		wait for Clk_period;
		Addr <=  "0001101001001";
		Trees_din <= x"1800611c";
		wait for Clk_period;
		Addr <=  "0001101001010";
		Trees_din <= x"03fdd20c";
		wait for Clk_period;
		Addr <=  "0001101001011";
		Trees_din <= x"02fa7204";
		wait for Clk_period;
		Addr <=  "0001101001100";
		Trees_din <= x"ff6e0e0d";
		wait for Clk_period;
		Addr <=  "0001101001101";
		Trees_din <= x"07013e04";
		wait for Clk_period;
		Addr <=  "0001101001110";
		Trees_din <= x"fff50e0d";
		wait for Clk_period;
		Addr <=  "0001101001111";
		Trees_din <= x"00de0e0d";
		wait for Clk_period;
		Addr <=  "0001101010000";
		Trees_din <= x"05fe6808";
		wait for Clk_period;
		Addr <=  "0001101010001";
		Trees_din <= x"08003c04";
		wait for Clk_period;
		Addr <=  "0001101010010";
		Trees_din <= x"ff930e0d";
		wait for Clk_period;
		Addr <=  "0001101010011";
		Trees_din <= x"00fb0e0d";
		wait for Clk_period;
		Addr <=  "0001101010100";
		Trees_din <= x"1300b304";
		wait for Clk_period;
		Addr <=  "0001101010101";
		Trees_din <= x"00900e0d";
		wait for Clk_period;
		Addr <=  "0001101010110";
		Trees_din <= x"ffb50e0d";
		wait for Clk_period;
		Addr <=  "0001101010111";
		Trees_din <= x"09004a10";
		wait for Clk_period;
		Addr <=  "0001101011000";
		Trees_din <= x"02faef08";
		wait for Clk_period;
		Addr <=  "0001101011001";
		Trees_din <= x"04065604";
		wait for Clk_period;
		Addr <=  "0001101011010";
		Trees_din <= x"ff740e0d";
		wait for Clk_period;
		Addr <=  "0001101011011";
		Trees_din <= x"ffde0e0d";
		wait for Clk_period;
		Addr <=  "0001101011100";
		Trees_din <= x"02faf804";
		wait for Clk_period;
		Addr <=  "0001101011101";
		Trees_din <= x"01600e0d";
		wait for Clk_period;
		Addr <=  "0001101011110";
		Trees_din <= x"ffee0e0d";
		wait for Clk_period;
		Addr <=  "0001101011111";
		Trees_din <= x"06080c08";
		wait for Clk_period;
		Addr <=  "0001101100000";
		Trees_din <= x"1300b304";
		wait for Clk_period;
		Addr <=  "0001101100001";
		Trees_din <= x"012f0e0d";
		wait for Clk_period;
		Addr <=  "0001101100010";
		Trees_din <= x"ff990e0d";
		wait for Clk_period;
		Addr <=  "0001101100011";
		Trees_din <= x"08005204";
		wait for Clk_period;
		Addr <=  "0001101100100";
		Trees_din <= x"ff760e0d";
		wait for Clk_period;
		Addr <=  "0001101100101";
		Trees_din <= x"00910e0d";
		wait for Clk_period;
		Addr <=  "0001101100110";
		Trees_din <= x"00fe2420";
		wait for Clk_period;
		Addr <=  "0001101100111";
		Trees_din <= x"12004910";
		wait for Clk_period;
		Addr <=  "0001101101000";
		Trees_din <= x"01fd0b08";
		wait for Clk_period;
		Addr <=  "0001101101001";
		Trees_din <= x"16031a04";
		wait for Clk_period;
		Addr <=  "0001101101010";
		Trees_din <= x"ffc40e0d";
		wait for Clk_period;
		Addr <=  "0001101101011";
		Trees_din <= x"00cc0e0d";
		wait for Clk_period;
		Addr <=  "0001101101100";
		Trees_din <= x"03fc1b04";
		wait for Clk_period;
		Addr <=  "0001101101101";
		Trees_din <= x"00620e0d";
		wait for Clk_period;
		Addr <=  "0001101101110";
		Trees_din <= x"ffd70e0d";
		wait for Clk_period;
		Addr <=  "0001101101111";
		Trees_din <= x"02f99f08";
		wait for Clk_period;
		Addr <=  "0001101110000";
		Trees_din <= x"04051704";
		wait for Clk_period;
		Addr <=  "0001101110001";
		Trees_din <= x"00850e0d";
		wait for Clk_period;
		Addr <=  "0001101110010";
		Trees_din <= x"ffac0e0d";
		wait for Clk_period;
		Addr <=  "0001101110011";
		Trees_din <= x"13009e04";
		wait for Clk_period;
		Addr <=  "0001101110100";
		Trees_din <= x"00f20e0d";
		wait for Clk_period;
		Addr <=  "0001101110101";
		Trees_din <= x"004d0e0d";
		wait for Clk_period;
		Addr <=  "0001101110110";
		Trees_din <= x"0707270c";
		wait for Clk_period;
		Addr <=  "0001101110111";
		Trees_din <= x"1b028708";
		wait for Clk_period;
		Addr <=  "0001101111000";
		Trees_din <= x"0a000b04";
		wait for Clk_period;
		Addr <=  "0001101111001";
		Trees_din <= x"00550e0d";
		wait for Clk_period;
		Addr <=  "0001101111010";
		Trees_din <= x"00080e0d";
		wait for Clk_period;
		Addr <=  "0001101111011";
		Trees_din <= x"ff620e0d";
		wait for Clk_period;
		Addr <=  "0001101111100";
		Trees_din <= x"02f8fa08";
		wait for Clk_period;
		Addr <=  "0001101111101";
		Trees_din <= x"07094904";
		wait for Clk_period;
		Addr <=  "0001101111110";
		Trees_din <= x"ffad0e0d";
		wait for Clk_period;
		Addr <=  "0001101111111";
		Trees_din <= x"006d0e0d";
		wait for Clk_period;
		Addr <=  "0001110000000";
		Trees_din <= x"0b00d704";
		wait for Clk_period;
		Addr <=  "0001110000001";
		Trees_din <= x"00a20e0d";
		wait for Clk_period;
		Addr <=  "0001110000010";
		Trees_din <= x"003d0e0d";
		wait for Clk_period;
		Addr <=  "0001110000011";
		Trees_din <= x"07ff5540";
		wait for Clk_period;
		Addr <=  "0001110000100";
		Trees_din <= x"07fcd514";
		wait for Clk_period;
		Addr <=  "0001110000101";
		Trees_din <= x"1c02410c";
		wait for Clk_period;
		Addr <=  "0001110000110";
		Trees_din <= x"06066c08";
		wait for Clk_period;
		Addr <=  "0001110000111";
		Trees_din <= x"06032c04";
		wait for Clk_period;
		Addr <=  "0001110001000";
		Trees_din <= x"000e0f41";
		wait for Clk_period;
		Addr <=  "0001110001001";
		Trees_din <= x"00ae0f41";
		wait for Clk_period;
		Addr <=  "0001110001010";
		Trees_din <= x"ff940f41";
		wait for Clk_period;
		Addr <=  "0001110001011";
		Trees_din <= x"12003004";
		wait for Clk_period;
		Addr <=  "0001110001100";
		Trees_din <= x"00430f41";
		wait for Clk_period;
		Addr <=  "0001110001101";
		Trees_din <= x"ff690f41";
		wait for Clk_period;
		Addr <=  "0001110001110";
		Trees_din <= x"1c026214";
		wait for Clk_period;
		Addr <=  "0001110001111";
		Trees_din <= x"0406840c";
		wait for Clk_period;
		Addr <=  "0001110010000";
		Trees_din <= x"0a016304";
		wait for Clk_period;
		Addr <=  "0001110010001";
		Trees_din <= x"ff680f41";
		wait for Clk_period;
		Addr <=  "0001110010010";
		Trees_din <= x"00fd4404";
		wait for Clk_period;
		Addr <=  "0001110010011";
		Trees_din <= x"00400f41";
		wait for Clk_period;
		Addr <=  "0001110010100";
		Trees_din <= x"ff950f41";
		wait for Clk_period;
		Addr <=  "0001110010101";
		Trees_din <= x"11000004";
		wait for Clk_period;
		Addr <=  "0001110010110";
		Trees_din <= x"00c90f41";
		wait for Clk_period;
		Addr <=  "0001110010111";
		Trees_din <= x"ff8d0f41";
		wait for Clk_period;
		Addr <=  "0001110011000";
		Trees_din <= x"1c026408";
		wait for Clk_period;
		Addr <=  "0001110011001";
		Trees_din <= x"04039304";
		wait for Clk_period;
		Addr <=  "0001110011010";
		Trees_din <= x"006d0f41";
		wait for Clk_period;
		Addr <=  "0001110011011";
		Trees_din <= x"01e60f41";
		wait for Clk_period;
		Addr <=  "0001110011100";
		Trees_din <= x"12004708";
		wait for Clk_period;
		Addr <=  "0001110011101";
		Trees_din <= x"00fc5604";
		wait for Clk_period;
		Addr <=  "0001110011110";
		Trees_din <= x"01220f41";
		wait for Clk_period;
		Addr <=  "0001110011111";
		Trees_din <= x"ff930f41";
		wait for Clk_period;
		Addr <=  "0001110100000";
		Trees_din <= x"18006a04";
		wait for Clk_period;
		Addr <=  "0001110100001";
		Trees_din <= x"01170f41";
		wait for Clk_period;
		Addr <=  "0001110100010";
		Trees_din <= x"ffff0f41";
		wait for Clk_period;
		Addr <=  "0001110100011";
		Trees_din <= x"0707273c";
		wait for Clk_period;
		Addr <=  "0001110100100";
		Trees_din <= x"02faca1c";
		wait for Clk_period;
		Addr <=  "0001110100101";
		Trees_din <= x"0e004510";
		wait for Clk_period;
		Addr <=  "0001110100110";
		Trees_din <= x"0e002108";
		wait for Clk_period;
		Addr <=  "0001110100111";
		Trees_din <= x"0e002104";
		wait for Clk_period;
		Addr <=  "0001110101000";
		Trees_din <= x"002d0f41";
		wait for Clk_period;
		Addr <=  "0001110101001";
		Trees_din <= x"01530f41";
		wait for Clk_period;
		Addr <=  "0001110101010";
		Trees_din <= x"16038904";
		wait for Clk_period;
		Addr <=  "0001110101011";
		Trees_din <= x"00260f41";
		wait for Clk_period;
		Addr <=  "0001110101100";
		Trees_din <= x"ffcb0f41";
		wait for Clk_period;
		Addr <=  "0001110101101";
		Trees_din <= x"0f007108";
		wait for Clk_period;
		Addr <=  "0001110101110";
		Trees_din <= x"0701d104";
		wait for Clk_period;
		Addr <=  "0001110101111";
		Trees_din <= x"ffa10f41";
		wait for Clk_period;
		Addr <=  "0001110110000";
		Trees_din <= x"00700f41";
		wait for Clk_period;
		Addr <=  "0001110110001";
		Trees_din <= x"01390f41";
		wait for Clk_period;
		Addr <=  "0001110110010";
		Trees_din <= x"19000e10";
		wait for Clk_period;
		Addr <=  "0001110110011";
		Trees_din <= x"060a9908";
		wait for Clk_period;
		Addr <=  "0001110110100";
		Trees_din <= x"1c022f04";
		wait for Clk_period;
		Addr <=  "0001110110101";
		Trees_din <= x"ff760f41";
		wait for Clk_period;
		Addr <=  "0001110110110";
		Trees_din <= x"00420f41";
		wait for Clk_period;
		Addr <=  "0001110110111";
		Trees_din <= x"08003b04";
		wait for Clk_period;
		Addr <=  "0001110111000";
		Trees_din <= x"01240f41";
		wait for Clk_period;
		Addr <=  "0001110111001";
		Trees_din <= x"ff910f41";
		wait for Clk_period;
		Addr <=  "0001110111010";
		Trees_din <= x"07021908";
		wait for Clk_period;
		Addr <=  "0001110111011";
		Trees_din <= x"1f028804";
		wait for Clk_period;
		Addr <=  "0001110111100";
		Trees_din <= x"ff7b0f41";
		wait for Clk_period;
		Addr <=  "0001110111101";
		Trees_din <= x"00a50f41";
		wait for Clk_period;
		Addr <=  "0001110111110";
		Trees_din <= x"01fde104";
		wait for Clk_period;
		Addr <=  "0001110111111";
		Trees_din <= x"006a0f41";
		wait for Clk_period;
		Addr <=  "0001111000000";
		Trees_din <= x"ffc90f41";
		wait for Clk_period;
		Addr <=  "0001111000001";
		Trees_din <= x"20040008";
		wait for Clk_period;
		Addr <=  "0001111000010";
		Trees_din <= x"0402d004";
		wait for Clk_period;
		Addr <=  "0001111000011";
		Trees_din <= x"003a0f41";
		wait for Clk_period;
		Addr <=  "0001111000100";
		Trees_din <= x"00b30f41";
		wait for Clk_period;
		Addr <=  "0001111000101";
		Trees_din <= x"02f8bf08";
		wait for Clk_period;
		Addr <=  "0001111000110";
		Trees_din <= x"07094904";
		wait for Clk_period;
		Addr <=  "0001111000111";
		Trees_din <= x"ff390f41";
		wait for Clk_period;
		Addr <=  "0001111001000";
		Trees_din <= x"005e0f41";
		wait for Clk_period;
		Addr <=  "0001111001001";
		Trees_din <= x"01ff5908";
		wait for Clk_period;
		Addr <=  "0001111001010";
		Trees_din <= x"05fbbf04";
		wait for Clk_period;
		Addr <=  "0001111001011";
		Trees_din <= x"fffc0f41";
		wait for Clk_period;
		Addr <=  "0001111001100";
		Trees_din <= x"00aa0f41";
		wait for Clk_period;
		Addr <=  "0001111001101";
		Trees_din <= x"01ffbf04";
		wait for Clk_period;
		Addr <=  "0001111001110";
		Trees_din <= x"ff8e0f41";
		wait for Clk_period;
		Addr <=  "0001111001111";
		Trees_din <= x"004b0f41";
		wait for Clk_period;
		Addr <=  "0001111010000";
		Trees_din <= x"07fdaa1c";
		wait for Clk_period;
		Addr <=  "0001111010001";
		Trees_din <= x"0f007a04";
		wait for Clk_period;
		Addr <=  "0001111010010";
		Trees_din <= x"ff6b1055";
		wait for Clk_period;
		Addr <=  "0001111010011";
		Trees_din <= x"03054208";
		wait for Clk_period;
		Addr <=  "0001111010100";
		Trees_din <= x"0b00e304";
		wait for Clk_period;
		Addr <=  "0001111010101";
		Trees_din <= x"ff741055";
		wait for Clk_period;
		Addr <=  "0001111010110";
		Trees_din <= x"00391055";
		wait for Clk_period;
		Addr <=  "0001111010111";
		Trees_din <= x"07fa6604";
		wait for Clk_period;
		Addr <=  "0001111011000";
		Trees_din <= x"ff8c1055";
		wait for Clk_period;
		Addr <=  "0001111011001";
		Trees_din <= x"0a016008";
		wait for Clk_period;
		Addr <=  "0001111011010";
		Trees_din <= x"1c024004";
		wait for Clk_period;
		Addr <=  "0001111011011";
		Trees_din <= x"00931055";
		wait for Clk_period;
		Addr <=  "0001111011100";
		Trees_din <= x"ffa11055";
		wait for Clk_period;
		Addr <=  "0001111011101";
		Trees_din <= x"012a1055";
		wait for Clk_period;
		Addr <=  "0001111011110";
		Trees_din <= x"07018e38";
		wait for Clk_period;
		Addr <=  "0001111011111";
		Trees_din <= x"03fbe918";
		wait for Clk_period;
		Addr <=  "0001111100000";
		Trees_din <= x"0c020a0c";
		wait for Clk_period;
		Addr <=  "0001111100001";
		Trees_din <= x"1d028808";
		wait for Clk_period;
		Addr <=  "0001111100010";
		Trees_din <= x"05fce504";
		wait for Clk_period;
		Addr <=  "0001111100011";
		Trees_din <= x"ffd91055";
		wait for Clk_period;
		Addr <=  "0001111100100";
		Trees_din <= x"ff611055";
		wait for Clk_period;
		Addr <=  "0001111100101";
		Trees_din <= x"00ad1055";
		wait for Clk_period;
		Addr <=  "0001111100110";
		Trees_din <= x"06090c08";
		wait for Clk_period;
		Addr <=  "0001111100111";
		Trees_din <= x"0406be04";
		wait for Clk_period;
		Addr <=  "0001111101000";
		Trees_din <= x"00ed1055";
		wait for Clk_period;
		Addr <=  "0001111101001";
		Trees_din <= x"ffe61055";
		wait for Clk_period;
		Addr <=  "0001111101010";
		Trees_din <= x"ff7b1055";
		wait for Clk_period;
		Addr <=  "0001111101011";
		Trees_din <= x"09004a10";
		wait for Clk_period;
		Addr <=  "0001111101100";
		Trees_din <= x"02fa5c08";
		wait for Clk_period;
		Addr <=  "0001111101101";
		Trees_din <= x"19005404";
		wait for Clk_period;
		Addr <=  "0001111101110";
		Trees_din <= x"ff801055";
		wait for Clk_period;
		Addr <=  "0001111101111";
		Trees_din <= x"00d41055";
		wait for Clk_period;
		Addr <=  "0001111110000";
		Trees_din <= x"0f005b04";
		wait for Clk_period;
		Addr <=  "0001111110001";
		Trees_din <= x"00b11055";
		wait for Clk_period;
		Addr <=  "0001111110010";
		Trees_din <= x"00051055";
		wait for Clk_period;
		Addr <=  "0001111110011";
		Trees_din <= x"00ff1808";
		wait for Clk_period;
		Addr <=  "0001111110100";
		Trees_din <= x"13009504";
		wait for Clk_period;
		Addr <=  "0001111110101";
		Trees_din <= x"ff9b1055";
		wait for Clk_period;
		Addr <=  "0001111110110";
		Trees_din <= x"00d91055";
		wait for Clk_period;
		Addr <=  "0001111110111";
		Trees_din <= x"22000804";
		wait for Clk_period;
		Addr <=  "0001111111000";
		Trees_din <= x"ff791055";
		wait for Clk_period;
		Addr <=  "0001111111001";
		Trees_din <= x"00801055";
		wait for Clk_period;
		Addr <=  "0001111111010";
		Trees_din <= x"00fe2418";
		wait for Clk_period;
		Addr <=  "0001111111011";
		Trees_din <= x"02f8fa08";
		wait for Clk_period;
		Addr <=  "0001111111100";
		Trees_din <= x"0b00d904";
		wait for Clk_period;
		Addr <=  "0001111111101";
		Trees_din <= x"ff661055";
		wait for Clk_period;
		Addr <=  "0001111111110";
		Trees_din <= x"002a1055";
		wait for Clk_period;
		Addr <=  "0001111111111";
		Trees_din <= x"1fff8708";
		wait for Clk_period;
		Addr <=  "0010000000000";
		Trees_din <= x"02fa9b04";
		wait for Clk_period;
		Addr <=  "0010000000001";
		Trees_din <= x"ff5c1055";
		wait for Clk_period;
		Addr <=  "0010000000010";
		Trees_din <= x"005d1055";
		wait for Clk_period;
		Addr <=  "0010000000011";
		Trees_din <= x"00fdf004";
		wait for Clk_period;
		Addr <=  "0010000000100";
		Trees_din <= x"004b1055";
		wait for Clk_period;
		Addr <=  "0010000000101";
		Trees_din <= x"00bb1055";
		wait for Clk_period;
		Addr <=  "0010000000110";
		Trees_din <= x"07072710";
		wait for Clk_period;
		Addr <=  "0010000000111";
		Trees_din <= x"05fe2b08";
		wait for Clk_period;
		Addr <=  "0010000001000";
		Trees_din <= x"06fca304";
		wait for Clk_period;
		Addr <=  "0010000001001";
		Trees_din <= x"ff8d1055";
		wait for Clk_period;
		Addr <=  "0010000001010";
		Trees_din <= x"000c1055";
		wait for Clk_period;
		Addr <=  "0010000001011";
		Trees_din <= x"0c011604";
		wait for Clk_period;
		Addr <=  "0010000001100";
		Trees_din <= x"008d1055";
		wait for Clk_period;
		Addr <=  "0010000001101";
		Trees_din <= x"fff51055";
		wait for Clk_period;
		Addr <=  "0010000001110";
		Trees_din <= x"20040008";
		wait for Clk_period;
		Addr <=  "0010000001111";
		Trees_din <= x"0402d004";
		wait for Clk_period;
		Addr <=  "0010000010000";
		Trees_din <= x"00321055";
		wait for Clk_period;
		Addr <=  "0010000010001";
		Trees_din <= x"00a91055";
		wait for Clk_period;
		Addr <=  "0010000010010";
		Trees_din <= x"08003f04";
		wait for Clk_period;
		Addr <=  "0010000010011";
		Trees_din <= x"00911055";
		wait for Clk_period;
		Addr <=  "0010000010100";
		Trees_din <= x"00191055";
		wait for Clk_period;
		Addr <=  "0010000010101";
		Trees_din <= x"07fdaa1c";
		wait for Clk_period;
		Addr <=  "0010000010110";
		Trees_din <= x"1800550c";
		wait for Clk_period;
		Addr <=  "0010000010111";
		Trees_din <= x"0d007c04";
		wait for Clk_period;
		Addr <=  "0010000011000";
		Trees_din <= x"00cc1151";
		wait for Clk_period;
		Addr <=  "0010000011001";
		Trees_din <= x"01fcbc04";
		wait for Clk_period;
		Addr <=  "0010000011010";
		Trees_din <= x"00421151";
		wait for Clk_period;
		Addr <=  "0010000011011";
		Trees_din <= x"ff831151";
		wait for Clk_period;
		Addr <=  "0010000011100";
		Trees_din <= x"04e87808";
		wait for Clk_period;
		Addr <=  "0010000011101";
		Trees_din <= x"07fbdc04";
		wait for Clk_period;
		Addr <=  "0010000011110";
		Trees_din <= x"ffa31151";
		wait for Clk_period;
		Addr <=  "0010000011111";
		Trees_din <= x"00841151";
		wait for Clk_period;
		Addr <=  "0010000100000";
		Trees_din <= x"0002d504";
		wait for Clk_period;
		Addr <=  "0010000100001";
		Trees_din <= x"ff6b1151";
		wait for Clk_period;
		Addr <=  "0010000100010";
		Trees_din <= x"00301151";
		wait for Clk_period;
		Addr <=  "0010000100011";
		Trees_din <= x"07037224";
		wait for Clk_period;
		Addr <=  "0010000100100";
		Trees_din <= x"03fae010";
		wait for Clk_period;
		Addr <=  "0010000100101";
		Trees_din <= x"1f027004";
		wait for Clk_period;
		Addr <=  "0010000100110";
		Trees_din <= x"ff641151";
		wait for Clk_period;
		Addr <=  "0010000100111";
		Trees_din <= x"1f027304";
		wait for Clk_period;
		Addr <=  "0010000101000";
		Trees_din <= x"00e11151";
		wait for Clk_period;
		Addr <=  "0010000101001";
		Trees_din <= x"05fe1f04";
		wait for Clk_period;
		Addr <=  "0010000101010";
		Trees_din <= x"ffa61151";
		wait for Clk_period;
		Addr <=  "0010000101011";
		Trees_din <= x"00981151";
		wait for Clk_period;
		Addr <=  "0010000101100";
		Trees_din <= x"02f93708";
		wait for Clk_period;
		Addr <=  "0010000101101";
		Trees_din <= x"0402dd04";
		wait for Clk_period;
		Addr <=  "0010000101110";
		Trees_din <= x"00081151";
		wait for Clk_period;
		Addr <=  "0010000101111";
		Trees_din <= x"ff571151";
		wait for Clk_period;
		Addr <=  "0010000110000";
		Trees_din <= x"060cd708";
		wait for Clk_period;
		Addr <=  "0010000110001";
		Trees_din <= x"08004004";
		wait for Clk_period;
		Addr <=  "0010000110010";
		Trees_din <= x"fff31151";
		wait for Clk_period;
		Addr <=  "0010000110011";
		Trees_din <= x"00201151";
		wait for Clk_period;
		Addr <=  "0010000110100";
		Trees_din <= x"ff791151";
		wait for Clk_period;
		Addr <=  "0010000110101";
		Trees_din <= x"19000120";
		wait for Clk_period;
		Addr <=  "0010000110110";
		Trees_din <= x"06019110";
		wait for Clk_period;
		Addr <=  "0010000110111";
		Trees_din <= x"15f81708";
		wait for Clk_period;
		Addr <=  "0010000111000";
		Trees_din <= x"0e002104";
		wait for Clk_period;
		Addr <=  "0010000111001";
		Trees_din <= x"00991151";
		wait for Clk_period;
		Addr <=  "0010000111010";
		Trees_din <= x"ffe81151";
		wait for Clk_period;
		Addr <=  "0010000111011";
		Trees_din <= x"14003104";
		wait for Clk_period;
		Addr <=  "0010000111100";
		Trees_din <= x"ffdf1151";
		wait for Clk_period;
		Addr <=  "0010000111101";
		Trees_din <= x"00941151";
		wait for Clk_period;
		Addr <=  "0010000111110";
		Trees_din <= x"01fcdf08";
		wait for Clk_period;
		Addr <=  "0010000111111";
		Trees_din <= x"1300a504";
		wait for Clk_period;
		Addr <=  "0010001000000";
		Trees_din <= x"00521151";
		wait for Clk_period;
		Addr <=  "0010001000001";
		Trees_din <= x"ff991151";
		wait for Clk_period;
		Addr <=  "0010001000010";
		Trees_din <= x"09002a04";
		wait for Clk_period;
		Addr <=  "0010001000011";
		Trees_din <= x"ff971151";
		wait for Clk_period;
		Addr <=  "0010001000100";
		Trees_din <= x"00b71151";
		wait for Clk_period;
		Addr <=  "0010001000101";
		Trees_din <= x"09004510";
		wait for Clk_period;
		Addr <=  "0010001000110";
		Trees_din <= x"1603f608";
		wait for Clk_period;
		Addr <=  "0010001000111";
		Trees_din <= x"02fb5f04";
		wait for Clk_period;
		Addr <=  "0010001001000";
		Trees_din <= x"00701151";
		wait for Clk_period;
		Addr <=  "0010001001001";
		Trees_din <= x"ffbf1151";
		wait for Clk_period;
		Addr <=  "0010001001010";
		Trees_din <= x"13009f04";
		wait for Clk_period;
		Addr <=  "0010001001011";
		Trees_din <= x"00961151";
		wait for Clk_period;
		Addr <=  "0010001001100";
		Trees_din <= x"ff8a1151";
		wait for Clk_period;
		Addr <=  "0010001001101";
		Trees_din <= x"00013608";
		wait for Clk_period;
		Addr <=  "0010001001110";
		Trees_din <= x"0a024504";
		wait for Clk_period;
		Addr <=  "0010001001111";
		Trees_din <= x"ff3a1151";
		wait for Clk_period;
		Addr <=  "0010001010000";
		Trees_din <= x"ffe91151";
		wait for Clk_period;
		Addr <=  "0010001010001";
		Trees_din <= x"05fd3a04";
		wait for Clk_period;
		Addr <=  "0010001010010";
		Trees_din <= x"ffa71151";
		wait for Clk_period;
		Addr <=  "0010001010011";
		Trees_din <= x"00781151";
		wait for Clk_period;
		Addr <=  "0010001010100";
		Trees_din <= x"07fdaa1c";
		wait for Clk_period;
		Addr <=  "0010001010101";
		Trees_din <= x"0f007a04";
		wait for Clk_period;
		Addr <=  "0010001010110";
		Trees_din <= x"ff6e1265";
		wait for Clk_period;
		Addr <=  "0010001010111";
		Trees_din <= x"03054208";
		wait for Clk_period;
		Addr <=  "0010001011000";
		Trees_din <= x"0b00e304";
		wait for Clk_period;
		Addr <=  "0010001011001";
		Trees_din <= x"ff7a1265";
		wait for Clk_period;
		Addr <=  "0010001011010";
		Trees_din <= x"00371265";
		wait for Clk_period;
		Addr <=  "0010001011011";
		Trees_din <= x"07fa6604";
		wait for Clk_period;
		Addr <=  "0010001011100";
		Trees_din <= x"ff981265";
		wait for Clk_period;
		Addr <=  "0010001011101";
		Trees_din <= x"0a016008";
		wait for Clk_period;
		Addr <=  "0010001011110";
		Trees_din <= x"1c024004";
		wait for Clk_period;
		Addr <=  "0010001011111";
		Trees_din <= x"00761265";
		wait for Clk_period;
		Addr <=  "0010001100000";
		Trees_din <= x"ffad1265";
		wait for Clk_period;
		Addr <=  "0010001100001";
		Trees_din <= x"00ea1265";
		wait for Clk_period;
		Addr <=  "0010001100010";
		Trees_din <= x"0e00213c";
		wait for Clk_period;
		Addr <=  "0010001100011";
		Trees_din <= x"00fe8120";
		wait for Clk_period;
		Addr <=  "0010001100100";
		Trees_din <= x"00fdfd10";
		wait for Clk_period;
		Addr <=  "0010001100101";
		Trees_din <= x"06050908";
		wait for Clk_period;
		Addr <=  "0010001100110";
		Trees_din <= x"1b027404";
		wait for Clk_period;
		Addr <=  "0010001100111";
		Trees_din <= x"00c01265";
		wait for Clk_period;
		Addr <=  "0010001101000";
		Trees_din <= x"ffbe1265";
		wait for Clk_period;
		Addr <=  "0010001101001";
		Trees_din <= x"12003804";
		wait for Clk_period;
		Addr <=  "0010001101010";
		Trees_din <= x"ff691265";
		wait for Clk_period;
		Addr <=  "0010001101011";
		Trees_din <= x"003f1265";
		wait for Clk_period;
		Addr <=  "0010001101100";
		Trees_din <= x"10002408";
		wait for Clk_period;
		Addr <=  "0010001101101";
		Trees_din <= x"15f72504";
		wait for Clk_period;
		Addr <=  "0010001101110";
		Trees_din <= x"00ba1265";
		wait for Clk_period;
		Addr <=  "0010001101111";
		Trees_din <= x"ffa31265";
		wait for Clk_period;
		Addr <=  "0010001110000";
		Trees_din <= x"1702ff04";
		wait for Clk_period;
		Addr <=  "0010001110001";
		Trees_din <= x"00031265";
		wait for Clk_period;
		Addr <=  "0010001110010";
		Trees_din <= x"014b1265";
		wait for Clk_period;
		Addr <=  "0010001110011";
		Trees_din <= x"0d009d10";
		wait for Clk_period;
		Addr <=  "0010001110100";
		Trees_din <= x"0b00d408";
		wait for Clk_period;
		Addr <=  "0010001110101";
		Trees_din <= x"08004204";
		wait for Clk_period;
		Addr <=  "0010001110110";
		Trees_din <= x"ffd81265";
		wait for Clk_period;
		Addr <=  "0010001110111";
		Trees_din <= x"00d01265";
		wait for Clk_period;
		Addr <=  "0010001111000";
		Trees_din <= x"0703f704";
		wait for Clk_period;
		Addr <=  "0010001111001";
		Trees_din <= x"ffc31265";
		wait for Clk_period;
		Addr <=  "0010001111010";
		Trees_din <= x"006d1265";
		wait for Clk_period;
		Addr <=  "0010001111011";
		Trees_din <= x"1002a608";
		wait for Clk_period;
		Addr <=  "0010001111100";
		Trees_din <= x"16040004";
		wait for Clk_period;
		Addr <=  "0010001111101";
		Trees_din <= x"ff741265";
		wait for Clk_period;
		Addr <=  "0010001111110";
		Trees_din <= x"00191265";
		wait for Clk_period;
		Addr <=  "0010001111111";
		Trees_din <= x"00481265";
		wait for Clk_period;
		Addr <=  "0010010000000";
		Trees_din <= x"2003fe14";
		wait for Clk_period;
		Addr <=  "0010010000001";
		Trees_din <= x"22004c08";
		wait for Clk_period;
		Addr <=  "0010010000010";
		Trees_din <= x"10004204";
		wait for Clk_period;
		Addr <=  "0010010000011";
		Trees_din <= x"01861265";
		wait for Clk_period;
		Addr <=  "0010010000100";
		Trees_din <= x"00741265";
		wait for Clk_period;
		Addr <=  "0010010000101";
		Trees_din <= x"1300b008";
		wait for Clk_period;
		Addr <=  "0010010000110";
		Trees_din <= x"09004a04";
		wait for Clk_period;
		Addr <=  "0010010000111";
		Trees_din <= x"00bc1265";
		wait for Clk_period;
		Addr <=  "0010010001000";
		Trees_din <= x"00061265";
		wait for Clk_period;
		Addr <=  "0010010001001";
		Trees_din <= x"ff671265";
		wait for Clk_period;
		Addr <=  "0010010001010";
		Trees_din <= x"07072710";
		wait for Clk_period;
		Addr <=  "0010010001011";
		Trees_din <= x"00fd3d08";
		wait for Clk_period;
		Addr <=  "0010010001100";
		Trees_din <= x"09003904";
		wait for Clk_period;
		Addr <=  "0010010001101";
		Trees_din <= x"ffb71265";
		wait for Clk_period;
		Addr <=  "0010010001110";
		Trees_din <= x"004d1265";
		wait for Clk_period;
		Addr <=  "0010010001111";
		Trees_din <= x"0b009404";
		wait for Clk_period;
		Addr <=  "0010010010000";
		Trees_din <= x"ffc91265";
		wait for Clk_period;
		Addr <=  "0010010010001";
		Trees_din <= x"00041265";
		wait for Clk_period;
		Addr <=  "0010010010010";
		Trees_din <= x"02f8fa08";
		wait for Clk_period;
		Addr <=  "0010010010011";
		Trees_din <= x"08004204";
		wait for Clk_period;
		Addr <=  "0010010010100";
		Trees_din <= x"00701265";
		wait for Clk_period;
		Addr <=  "0010010010101";
		Trees_din <= x"ffa11265";
		wait for Clk_period;
		Addr <=  "0010010010110";
		Trees_din <= x"05fbbf04";
		wait for Clk_period;
		Addr <=  "0010010010111";
		Trees_din <= x"001c1265";
		wait for Clk_period;
		Addr <=  "0010010011000";
		Trees_din <= x"00811265";
		wait for Clk_period;
		Addr <=  "0010010011001";
		Trees_din <= x"07fcd510";
		wait for Clk_period;
		Addr <=  "0010010011010";
		Trees_din <= x"1300e608";
		wait for Clk_period;
		Addr <=  "0010010011011";
		Trees_din <= x"05157904";
		wait for Clk_period;
		Addr <=  "0010010011100";
		Trees_din <= x"ff6f1381";
		wait for Clk_period;
		Addr <=  "0010010011101";
		Trees_din <= x"00111381";
		wait for Clk_period;
		Addr <=  "0010010011110";
		Trees_din <= x"1300ea04";
		wait for Clk_period;
		Addr <=  "0010010011111";
		Trees_din <= x"009b1381";
		wait for Clk_period;
		Addr <=  "0010010100000";
		Trees_din <= x"ffb01381";
		wait for Clk_period;
		Addr <=  "0010010100001";
		Trees_din <= x"1d026b40";
		wait for Clk_period;
		Addr <=  "0010010100010";
		Trees_din <= x"1b026520";
		wait for Clk_period;
		Addr <=  "0010010100011";
		Trees_din <= x"03fb9310";
		wait for Clk_period;
		Addr <=  "0010010100100";
		Trees_din <= x"07021908";
		wait for Clk_period;
		Addr <=  "0010010100101";
		Trees_din <= x"0b00fe04";
		wait for Clk_period;
		Addr <=  "0010010100110";
		Trees_din <= x"ff651381";
		wait for Clk_period;
		Addr <=  "0010010100111";
		Trees_din <= x"00131381";
		wait for Clk_period;
		Addr <=  "0010010101000";
		Trees_din <= x"00ff3804";
		wait for Clk_period;
		Addr <=  "0010010101001";
		Trees_din <= x"00781381";
		wait for Clk_period;
		Addr <=  "0010010101010";
		Trees_din <= x"ffb11381";
		wait for Clk_period;
		Addr <=  "0010010101011";
		Trees_din <= x"01fc9c08";
		wait for Clk_period;
		Addr <=  "0010010101100";
		Trees_din <= x"0d007a04";
		wait for Clk_period;
		Addr <=  "0010010101101";
		Trees_din <= x"ff9a1381";
		wait for Clk_period;
		Addr <=  "0010010101110";
		Trees_din <= x"00491381";
		wait for Clk_period;
		Addr <=  "0010010101111";
		Trees_din <= x"1e026304";
		wait for Clk_period;
		Addr <=  "0010010110000";
		Trees_din <= x"00181381";
		wait for Clk_period;
		Addr <=  "0010010110001";
		Trees_din <= x"00711381";
		wait for Clk_period;
		Addr <=  "0010010110010";
		Trees_din <= x"00005010";
		wait for Clk_period;
		Addr <=  "0010010110011";
		Trees_din <= x"05fc5208";
		wait for Clk_period;
		Addr <=  "0010010110100";
		Trees_din <= x"1f026804";
		wait for Clk_period;
		Addr <=  "0010010110101";
		Trees_din <= x"ff9f1381";
		wait for Clk_period;
		Addr <=  "0010010110110";
		Trees_din <= x"00881381";
		wait for Clk_period;
		Addr <=  "0010010110111";
		Trees_din <= x"08005104";
		wait for Clk_period;
		Addr <=  "0010010111000";
		Trees_din <= x"ff6a1381";
		wait for Clk_period;
		Addr <=  "0010010111001";
		Trees_din <= x"fff01381";
		wait for Clk_period;
		Addr <=  "0010010111010";
		Trees_din <= x"0b00dc08";
		wait for Clk_period;
		Addr <=  "0010010111011";
		Trees_din <= x"12004f04";
		wait for Clk_period;
		Addr <=  "0010010111100";
		Trees_din <= x"00b81381";
		wait for Clk_period;
		Addr <=  "0010010111101";
		Trees_din <= x"ffcf1381";
		wait for Clk_period;
		Addr <=  "0010010111110";
		Trees_din <= x"05fd3e04";
		wait for Clk_period;
		Addr <=  "0010010111111";
		Trees_din <= x"ff821381";
		wait for Clk_period;
		Addr <=  "0010011000000";
		Trees_din <= x"004d1381";
		wait for Clk_period;
		Addr <=  "0010011000001";
		Trees_din <= x"0c012a20";
		wait for Clk_period;
		Addr <=  "0010011000010";
		Trees_din <= x"10007210";
		wait for Clk_period;
		Addr <=  "0010011000011";
		Trees_din <= x"1b027208";
		wait for Clk_period;
		Addr <=  "0010011000100";
		Trees_din <= x"0d007104";
		wait for Clk_period;
		Addr <=  "0010011000101";
		Trees_din <= x"ffb51381";
		wait for Clk_period;
		Addr <=  "0010011000110";
		Trees_din <= x"00911381";
		wait for Clk_period;
		Addr <=  "0010011000111";
		Trees_din <= x"09004c04";
		wait for Clk_period;
		Addr <=  "0010011001000";
		Trees_din <= x"ffbd1381";
		wait for Clk_period;
		Addr <=  "0010011001001";
		Trees_din <= x"00c31381";
		wait for Clk_period;
		Addr <=  "0010011001010";
		Trees_din <= x"10027008";
		wait for Clk_period;
		Addr <=  "0010011001011";
		Trees_din <= x"07017704";
		wait for Clk_period;
		Addr <=  "0010011001100";
		Trees_din <= x"004c1381";
		wait for Clk_period;
		Addr <=  "0010011001101";
		Trees_din <= x"00dc1381";
		wait for Clk_period;
		Addr <=  "0010011001110";
		Trees_din <= x"0e004404";
		wait for Clk_period;
		Addr <=  "0010011001111";
		Trees_din <= x"ffb61381";
		wait for Clk_period;
		Addr <=  "0010011010000";
		Trees_din <= x"00891381";
		wait for Clk_period;
		Addr <=  "0010011010001";
		Trees_din <= x"19000a10";
		wait for Clk_period;
		Addr <=  "0010011010010";
		Trees_din <= x"0c029608";
		wait for Clk_period;
		Addr <=  "0010011010011";
		Trees_din <= x"060b0c04";
		wait for Clk_period;
		Addr <=  "0010011010100";
		Trees_din <= x"00091381";
		wait for Clk_period;
		Addr <=  "0010011010101";
		Trees_din <= x"ff7a1381";
		wait for Clk_period;
		Addr <=  "0010011010110";
		Trees_din <= x"16038104";
		wait for Clk_period;
		Addr <=  "0010011010111";
		Trees_din <= x"00c41381";
		wait for Clk_period;
		Addr <=  "0010011011000";
		Trees_din <= x"001e1381";
		wait for Clk_period;
		Addr <=  "0010011011001";
		Trees_din <= x"18004f08";
		wait for Clk_period;
		Addr <=  "0010011011010";
		Trees_din <= x"1001b504";
		wait for Clk_period;
		Addr <=  "0010011011011";
		Trees_din <= x"00981381";
		wait for Clk_period;
		Addr <=  "0010011011100";
		Trees_din <= x"ffcf1381";
		wait for Clk_period;
		Addr <=  "0010011011101";
		Trees_din <= x"17029704";
		wait for Clk_period;
		Addr <=  "0010011011110";
		Trees_din <= x"000a1381";
		wait for Clk_period;
		Addr <=  "0010011011111";
		Trees_din <= x"ff831381";
		wait for Clk_period;
		Addr <=  "0010011100000";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0010011100001";
		Trees_din <= x"07fcd50c";
		wait for Clk_period;
		Addr <=  "0010011100010";
		Trees_din <= x"1300e608";
		wait for Clk_period;
		Addr <=  "0010011100011";
		Trees_din <= x"15f6f904";
		wait for Clk_period;
		Addr <=  "0010011100100";
		Trees_din <= x"001513f9";
		wait for Clk_period;
		Addr <=  "0010011100101";
		Trees_din <= x"ff7213f9";
		wait for Clk_period;
		Addr <=  "0010011100110";
		Trees_din <= x"002f13f9";
		wait for Clk_period;
		Addr <=  "0010011100111";
		Trees_din <= x"060cd72c";
		wait for Clk_period;
		Addr <=  "0010011101000";
		Trees_din <= x"15f6ca0c";
		wait for Clk_period;
		Addr <=  "0010011101001";
		Trees_din <= x"1f021004";
		wait for Clk_period;
		Addr <=  "0010011101010";
		Trees_din <= x"005913f9";
		wait for Clk_period;
		Addr <=  "0010011101011";
		Trees_din <= x"08004d04";
		wait for Clk_period;
		Addr <=  "0010011101100";
		Trees_din <= x"ff5f13f9";
		wait for Clk_period;
		Addr <=  "0010011101101";
		Trees_din <= x"000613f9";
		wait for Clk_period;
		Addr <=  "0010011101110";
		Trees_din <= x"15f6fc10";
		wait for Clk_period;
		Addr <=  "0010011101111";
		Trees_din <= x"01fd9908";
		wait for Clk_period;
		Addr <=  "0010011110000";
		Trees_din <= x"0e002804";
		wait for Clk_period;
		Addr <=  "0010011110001";
		Trees_din <= x"00c013f9";
		wait for Clk_period;
		Addr <=  "0010011110010";
		Trees_din <= x"ff7a13f9";
		wait for Clk_period;
		Addr <=  "0010011110011";
		Trees_din <= x"0b009704";
		wait for Clk_period;
		Addr <=  "0010011110100";
		Trees_din <= x"ff9f13f9";
		wait for Clk_period;
		Addr <=  "0010011110101";
		Trees_din <= x"00c013f9";
		wait for Clk_period;
		Addr <=  "0010011110110";
		Trees_din <= x"1d026b08";
		wait for Clk_period;
		Addr <=  "0010011110111";
		Trees_din <= x"0f007704";
		wait for Clk_period;
		Addr <=  "0010011111000";
		Trees_din <= x"ffdf13f9";
		wait for Clk_period;
		Addr <=  "0010011111001";
		Trees_din <= x"001513f9";
		wait for Clk_period;
		Addr <=  "0010011111010";
		Trees_din <= x"02fbce04";
		wait for Clk_period;
		Addr <=  "0010011111011";
		Trees_din <= x"000913f9";
		wait for Clk_period;
		Addr <=  "0010011111100";
		Trees_din <= x"004513f9";
		wait for Clk_period;
		Addr <=  "0010011111101";
		Trees_din <= x"ff7d13f9";
		wait for Clk_period;
		Addr <=  "0010011111110";
		Trees_din <= x"07018e64";
		wait for Clk_period;
		Addr <=  "0010011111111";
		Trees_din <= x"0a01ce40";
		wait for Clk_period;
		Addr <=  "0010100000000";
		Trees_din <= x"0a010920";
		wait for Clk_period;
		Addr <=  "0010100000001";
		Trees_din <= x"03fb9810";
		wait for Clk_period;
		Addr <=  "0010100000010";
		Trees_din <= x"17039408";
		wait for Clk_period;
		Addr <=  "0010100000011";
		Trees_din <= x"00fe4304";
		wait for Clk_period;
		Addr <=  "0010100000100";
		Trees_din <= x"00631565";
		wait for Clk_period;
		Addr <=  "0010100000101";
		Trees_din <= x"ff8f1565";
		wait for Clk_period;
		Addr <=  "0010100000110";
		Trees_din <= x"21000104";
		wait for Clk_period;
		Addr <=  "0010100000111";
		Trees_din <= x"ff671565";
		wait for Clk_period;
		Addr <=  "0010100001000";
		Trees_din <= x"00371565";
		wait for Clk_period;
		Addr <=  "0010100001001";
		Trees_din <= x"07fe4808";
		wait for Clk_period;
		Addr <=  "0010100001010";
		Trees_din <= x"0d007404";
		wait for Clk_period;
		Addr <=  "0010100001011";
		Trees_din <= x"ff701565";
		wait for Clk_period;
		Addr <=  "0010100001100";
		Trees_din <= x"ffec1565";
		wait for Clk_period;
		Addr <=  "0010100001101";
		Trees_din <= x"09003e04";
		wait for Clk_period;
		Addr <=  "0010100001110";
		Trees_din <= x"ffe71565";
		wait for Clk_period;
		Addr <=  "0010100001111";
		Trees_din <= x"00381565";
		wait for Clk_period;
		Addr <=  "0010100010000";
		Trees_din <= x"06070c10";
		wait for Clk_period;
		Addr <=  "0010100010001";
		Trees_din <= x"08004f08";
		wait for Clk_period;
		Addr <=  "0010100010010";
		Trees_din <= x"0000ee04";
		wait for Clk_period;
		Addr <=  "0010100010011";
		Trees_din <= x"ff781565";
		wait for Clk_period;
		Addr <=  "0010100010100";
		Trees_din <= x"004b1565";
		wait for Clk_period;
		Addr <=  "0010100010101";
		Trees_din <= x"0e003304";
		wait for Clk_period;
		Addr <=  "0010100010110";
		Trees_din <= x"00271565";
		wait for Clk_period;
		Addr <=  "0010100010111";
		Trees_din <= x"00c41565";
		wait for Clk_period;
		Addr <=  "0010100011000";
		Trees_din <= x"0a016008";
		wait for Clk_period;
		Addr <=  "0010100011001";
		Trees_din <= x"1d026204";
		wait for Clk_period;
		Addr <=  "0010100011010";
		Trees_din <= x"ffe31565";
		wait for Clk_period;
		Addr <=  "0010100011011";
		Trees_din <= x"01201565";
		wait for Clk_period;
		Addr <=  "0010100011100";
		Trees_din <= x"02fb8304";
		wait for Clk_period;
		Addr <=  "0010100011101";
		Trees_din <= x"ffa21565";
		wait for Clk_period;
		Addr <=  "0010100011110";
		Trees_din <= x"00881565";
		wait for Clk_period;
		Addr <=  "0010100011111";
		Trees_din <= x"1700c410";
		wait for Clk_period;
		Addr <=  "0010100100000";
		Trees_din <= x"02fbe308";
		wait for Clk_period;
		Addr <=  "0010100100001";
		Trees_din <= x"08004404";
		wait for Clk_period;
		Addr <=  "0010100100010";
		Trees_din <= x"002e1565";
		wait for Clk_period;
		Addr <=  "0010100100011";
		Trees_din <= x"ff871565";
		wait for Clk_period;
		Addr <=  "0010100100100";
		Trees_din <= x"1300b804";
		wait for Clk_period;
		Addr <=  "0010100100101";
		Trees_din <= x"01011565";
		wait for Clk_period;
		Addr <=  "0010100100110";
		Trees_din <= x"00251565";
		wait for Clk_period;
		Addr <=  "0010100100111";
		Trees_din <= x"1f028810";
		wait for Clk_period;
		Addr <=  "0010100101000";
		Trees_din <= x"09004b08";
		wait for Clk_period;
		Addr <=  "0010100101001";
		Trees_din <= x"0b00ab04";
		wait for Clk_period;
		Addr <=  "0010100101010";
		Trees_din <= x"ffbf1565";
		wait for Clk_period;
		Addr <=  "0010100101011";
		Trees_din <= x"ff621565";
		wait for Clk_period;
		Addr <=  "0010100101100";
		Trees_din <= x"0b007d04";
		wait for Clk_period;
		Addr <=  "0010100101101";
		Trees_din <= x"ff811565";
		wait for Clk_period;
		Addr <=  "0010100101110";
		Trees_din <= x"00a71565";
		wait for Clk_period;
		Addr <=  "0010100101111";
		Trees_din <= x"00951565";
		wait for Clk_period;
		Addr <=  "0010100110000";
		Trees_din <= x"0900342c";
		wait for Clk_period;
		Addr <=  "0010100110001";
		Trees_din <= x"18005c18";
		wait for Clk_period;
		Addr <=  "0010100110010";
		Trees_din <= x"0b00e710";
		wait for Clk_period;
		Addr <=  "0010100110011";
		Trees_din <= x"0d00a708";
		wait for Clk_period;
		Addr <=  "0010100110100";
		Trees_din <= x"07021904";
		wait for Clk_period;
		Addr <=  "0010100110101";
		Trees_din <= x"ffbb1565";
		wait for Clk_period;
		Addr <=  "0010100110110";
		Trees_din <= x"009d1565";
		wait for Clk_period;
		Addr <=  "0010100110111";
		Trees_din <= x"06ffea04";
		wait for Clk_period;
		Addr <=  "0010100111000";
		Trees_din <= x"00021565";
		wait for Clk_period;
		Addr <=  "0010100111001";
		Trees_din <= x"ff731565";
		wait for Clk_period;
		Addr <=  "0010100111010";
		Trees_din <= x"08004604";
		wait for Clk_period;
		Addr <=  "0010100111011";
		Trees_din <= x"ff5b1565";
		wait for Clk_period;
		Addr <=  "0010100111100";
		Trees_din <= x"00561565";
		wait for Clk_period;
		Addr <=  "0010100111101";
		Trees_din <= x"0701bc04";
		wait for Clk_period;
		Addr <=  "0010100111110";
		Trees_din <= x"ffcb1565";
		wait for Clk_period;
		Addr <=  "0010100111111";
		Trees_din <= x"0e002b08";
		wait for Clk_period;
		Addr <=  "0010101000000";
		Trees_din <= x"05fb7304";
		wait for Clk_period;
		Addr <=  "0010101000001";
		Trees_din <= x"ffc91565";
		wait for Clk_period;
		Addr <=  "0010101000010";
		Trees_din <= x"00bf1565";
		wait for Clk_period;
		Addr <=  "0010101000011";
		Trees_din <= x"13005b04";
		wait for Clk_period;
		Addr <=  "0010101000100";
		Trees_din <= x"00671565";
		wait for Clk_period;
		Addr <=  "0010101000101";
		Trees_din <= x"ffa21565";
		wait for Clk_period;
		Addr <=  "0010101000110";
		Trees_din <= x"1601290c";
		wait for Clk_period;
		Addr <=  "0010101000111";
		Trees_din <= x"1d002204";
		wait for Clk_period;
		Addr <=  "0010101001000";
		Trees_din <= x"ffdf1565";
		wait for Clk_period;
		Addr <=  "0010101001001";
		Trees_din <= x"01fe7904";
		wait for Clk_period;
		Addr <=  "0010101001010";
		Trees_din <= x"00e01565";
		wait for Clk_period;
		Addr <=  "0010101001011";
		Trees_din <= x"00041565";
		wait for Clk_period;
		Addr <=  "0010101001100";
		Trees_din <= x"15fa7f10";
		wait for Clk_period;
		Addr <=  "0010101001101";
		Trees_din <= x"0701aa08";
		wait for Clk_period;
		Addr <=  "0010101001110";
		Trees_din <= x"0a00fd04";
		wait for Clk_period;
		Addr <=  "0010101001111";
		Trees_din <= x"001a1565";
		wait for Clk_period;
		Addr <=  "0010101010000";
		Trees_din <= x"01261565";
		wait for Clk_period;
		Addr <=  "0010101010001";
		Trees_din <= x"09003904";
		wait for Clk_period;
		Addr <=  "0010101010010";
		Trees_din <= x"ffc11565";
		wait for Clk_period;
		Addr <=  "0010101010011";
		Trees_din <= x"00141565";
		wait for Clk_period;
		Addr <=  "0010101010100";
		Trees_din <= x"19000304";
		wait for Clk_period;
		Addr <=  "0010101010101";
		Trees_din <= x"00551565";
		wait for Clk_period;
		Addr <=  "0010101010110";
		Trees_din <= x"1300ae04";
		wait for Clk_period;
		Addr <=  "0010101010111";
		Trees_din <= x"00161565";
		wait for Clk_period;
		Addr <=  "0010101011000";
		Trees_din <= x"ff501565";
		wait for Clk_period;
		Addr <=  "0010101011001";
		Trees_din <= x"07fcd50c";
		wait for Clk_period;
		Addr <=  "0010101011010";
		Trees_din <= x"1300e608";
		wait for Clk_period;
		Addr <=  "0010101011011";
		Trees_din <= x"05157904";
		wait for Clk_period;
		Addr <=  "0010101011100";
		Trees_din <= x"ff751639";
		wait for Clk_period;
		Addr <=  "0010101011101";
		Trees_din <= x"001d1639";
		wait for Clk_period;
		Addr <=  "0010101011110";
		Trees_din <= x"002a1639";
		wait for Clk_period;
		Addr <=  "0010101011111";
		Trees_din <= x"0e002124";
		wait for Clk_period;
		Addr <=  "0010101100000";
		Trees_din <= x"0d007c04";
		wait for Clk_period;
		Addr <=  "0010101100001";
		Trees_din <= x"00fe1639";
		wait for Clk_period;
		Addr <=  "0010101100010";
		Trees_din <= x"08004210";
		wait for Clk_period;
		Addr <=  "0010101100011";
		Trees_din <= x"21000008";
		wait for Clk_period;
		Addr <=  "0010101100100";
		Trees_din <= x"16038d04";
		wait for Clk_period;
		Addr <=  "0010101100101";
		Trees_din <= x"ff7d1639";
		wait for Clk_period;
		Addr <=  "0010101100110";
		Trees_din <= x"fff51639";
		wait for Clk_period;
		Addr <=  "0010101100111";
		Trees_din <= x"0a000804";
		wait for Clk_period;
		Addr <=  "0010101101000";
		Trees_din <= x"00ce1639";
		wait for Clk_period;
		Addr <=  "0010101101001";
		Trees_din <= x"001b1639";
		wait for Clk_period;
		Addr <=  "0010101101010";
		Trees_din <= x"08004408";
		wait for Clk_period;
		Addr <=  "0010101101011";
		Trees_din <= x"11001404";
		wait for Clk_period;
		Addr <=  "0010101101100";
		Trees_din <= x"fffd1639";
		wait for Clk_period;
		Addr <=  "0010101101101";
		Trees_din <= x"00fd1639";
		wait for Clk_period;
		Addr <=  "0010101101110";
		Trees_din <= x"07015b04";
		wait for Clk_period;
		Addr <=  "0010101101111";
		Trees_din <= x"ffe21639";
		wait for Clk_period;
		Addr <=  "0010101110000";
		Trees_din <= x"004d1639";
		wait for Clk_period;
		Addr <=  "0010101110001";
		Trees_din <= x"1300be1c";
		wait for Clk_period;
		Addr <=  "0010101110010";
		Trees_din <= x"1400340c";
		wait for Clk_period;
		Addr <=  "0010101110011";
		Trees_din <= x"1300bd08";
		wait for Clk_period;
		Addr <=  "0010101110100";
		Trees_din <= x"19000604";
		wait for Clk_period;
		Addr <=  "0010101110101";
		Trees_din <= x"ff3e1639";
		wait for Clk_period;
		Addr <=  "0010101110110";
		Trees_din <= x"ffc51639";
		wait for Clk_period;
		Addr <=  "0010101110111";
		Trees_din <= x"007b1639";
		wait for Clk_period;
		Addr <=  "0010101111000";
		Trees_din <= x"14003808";
		wait for Clk_period;
		Addr <=  "0010101111001";
		Trees_din <= x"06075e04";
		wait for Clk_period;
		Addr <=  "0010101111010";
		Trees_din <= x"00961639";
		wait for Clk_period;
		Addr <=  "0010101111011";
		Trees_din <= x"ffe51639";
		wait for Clk_period;
		Addr <=  "0010101111100";
		Trees_din <= x"0b006304";
		wait for Clk_period;
		Addr <=  "0010101111101";
		Trees_din <= x"006b1639";
		wait for Clk_period;
		Addr <=  "0010101111110";
		Trees_din <= x"00021639";
		wait for Clk_period;
		Addr <=  "0010101111111";
		Trees_din <= x"12003910";
		wait for Clk_period;
		Addr <=  "0010110000000";
		Trees_din <= x"1703d908";
		wait for Clk_period;
		Addr <=  "0010110000001";
		Trees_din <= x"07016304";
		wait for Clk_period;
		Addr <=  "0010110000010";
		Trees_din <= x"ff7a1639";
		wait for Clk_period;
		Addr <=  "0010110000011";
		Trees_din <= x"004e1639";
		wait for Clk_period;
		Addr <=  "0010110000100";
		Trees_din <= x"08004004";
		wait for Clk_period;
		Addr <=  "0010110000101";
		Trees_din <= x"ffd81639";
		wait for Clk_period;
		Addr <=  "0010110000110";
		Trees_din <= x"01241639";
		wait for Clk_period;
		Addr <=  "0010110000111";
		Trees_din <= x"03031e08";
		wait for Clk_period;
		Addr <=  "0010110001000";
		Trees_din <= x"07072704";
		wait for Clk_period;
		Addr <=  "0010110001001";
		Trees_din <= x"ffa21639";
		wait for Clk_period;
		Addr <=  "0010110001010";
		Trees_din <= x"005b1639";
		wait for Clk_period;
		Addr <=  "0010110001011";
		Trees_din <= x"0606d104";
		wait for Clk_period;
		Addr <=  "0010110001100";
		Trees_din <= x"002b1639";
		wait for Clk_period;
		Addr <=  "0010110001101";
		Trees_din <= x"01381639";
		wait for Clk_period;
		Addr <=  "0010110001110";
		Trees_din <= x"07031054";
		wait for Clk_period;
		Addr <=  "0010110001111";
		Trees_din <= x"00ffd224";
		wait for Clk_period;
		Addr <=  "0010110010000";
		Trees_din <= x"07fdaa10";
		wait for Clk_period;
		Addr <=  "0010110010001";
		Trees_din <= x"00fc8f08";
		wait for Clk_period;
		Addr <=  "0010110010010";
		Trees_din <= x"0f008204";
		wait for Clk_period;
		Addr <=  "0010110010011";
		Trees_din <= x"ffa71795";
		wait for Clk_period;
		Addr <=  "0010110010100";
		Trees_din <= x"00861795";
		wait for Clk_period;
		Addr <=  "0010110010101";
		Trees_din <= x"1dff8204";
		wait for Clk_period;
		Addr <=  "0010110010110";
		Trees_din <= x"00041795";
		wait for Clk_period;
		Addr <=  "0010110010111";
		Trees_din <= x"ff741795";
		wait for Clk_period;
		Addr <=  "0010110011000";
		Trees_din <= x"02f91404";
		wait for Clk_period;
		Addr <=  "0010110011001";
		Trees_din <= x"ff6e1795";
		wait for Clk_period;
		Addr <=  "0010110011010";
		Trees_din <= x"00ff5c08";
		wait for Clk_period;
		Addr <=  "0010110011011";
		Trees_din <= x"09004904";
		wait for Clk_period;
		Addr <=  "0010110011100";
		Trees_din <= x"ffff1795";
		wait for Clk_period;
		Addr <=  "0010110011101";
		Trees_din <= x"004e1795";
		wait for Clk_period;
		Addr <=  "0010110011110";
		Trees_din <= x"05fdba04";
		wait for Clk_period;
		Addr <=  "0010110011111";
		Trees_din <= x"008d1795";
		wait for Clk_period;
		Addr <=  "0010110100000";
		Trees_din <= x"ffda1795";
		wait for Clk_period;
		Addr <=  "0010110100001";
		Trees_din <= x"00007210";
		wait for Clk_period;
		Addr <=  "0010110100010";
		Trees_din <= x"07ff7108";
		wait for Clk_period;
		Addr <=  "0010110100011";
		Trees_din <= x"0400fc04";
		wait for Clk_period;
		Addr <=  "0010110100100";
		Trees_din <= x"00921795";
		wait for Clk_period;
		Addr <=  "0010110100101";
		Trees_din <= x"ff931795";
		wait for Clk_period;
		Addr <=  "0010110100110";
		Trees_din <= x"03016c04";
		wait for Clk_period;
		Addr <=  "0010110100111";
		Trees_din <= x"ff571795";
		wait for Clk_period;
		Addr <=  "0010110101000";
		Trees_din <= x"ffe51795";
		wait for Clk_period;
		Addr <=  "0010110101001";
		Trees_din <= x"01fdec10";
		wait for Clk_period;
		Addr <=  "0010110101010";
		Trees_din <= x"0c01a108";
		wait for Clk_period;
		Addr <=  "0010110101011";
		Trees_din <= x"0c000404";
		wait for Clk_period;
		Addr <=  "0010110101100";
		Trees_din <= x"007b1795";
		wait for Clk_period;
		Addr <=  "0010110101101";
		Trees_din <= x"ff6f1795";
		wait for Clk_period;
		Addr <=  "0010110101110";
		Trees_din <= x"03fd4a04";
		wait for Clk_period;
		Addr <=  "0010110101111";
		Trees_din <= x"ffab1795";
		wait for Clk_period;
		Addr <=  "0010110110000";
		Trees_din <= x"00931795";
		wait for Clk_period;
		Addr <=  "0010110110001";
		Trees_din <= x"01fe5a08";
		wait for Clk_period;
		Addr <=  "0010110110010";
		Trees_din <= x"10000204";
		wait for Clk_period;
		Addr <=  "0010110110011";
		Trees_din <= x"ffe21795";
		wait for Clk_period;
		Addr <=  "0010110110100";
		Trees_din <= x"00ea1795";
		wait for Clk_period;
		Addr <=  "0010110110101";
		Trees_din <= x"05fd4204";
		wait for Clk_period;
		Addr <=  "0010110110110";
		Trees_din <= x"ff781795";
		wait for Clk_period;
		Addr <=  "0010110110111";
		Trees_din <= x"00181795";
		wait for Clk_period;
		Addr <=  "0010110111000";
		Trees_din <= x"0604c840";
		wait for Clk_period;
		Addr <=  "0010110111001";
		Trees_din <= x"1703d520";
		wait for Clk_period;
		Addr <=  "0010110111010";
		Trees_din <= x"1e025e10";
		wait for Clk_period;
		Addr <=  "0010110111011";
		Trees_din <= x"17031508";
		wait for Clk_period;
		Addr <=  "0010110111100";
		Trees_din <= x"04063804";
		wait for Clk_period;
		Addr <=  "0010110111101";
		Trees_din <= x"00501795";
		wait for Clk_period;
		Addr <=  "0010110111110";
		Trees_din <= x"ffb51795";
		wait for Clk_period;
		Addr <=  "0010110111111";
		Trees_din <= x"0c012504";
		wait for Clk_period;
		Addr <=  "0010111000000";
		Trees_din <= x"00431795";
		wait for Clk_period;
		Addr <=  "0010111000001";
		Trees_din <= x"00e21795";
		wait for Clk_period;
		Addr <=  "0010111000010";
		Trees_din <= x"19000108";
		wait for Clk_period;
		Addr <=  "0010111000011";
		Trees_din <= x"12004c04";
		wait for Clk_period;
		Addr <=  "0010111000100";
		Trees_din <= x"000a1795";
		wait for Clk_period;
		Addr <=  "0010111000101";
		Trees_din <= x"006c1795";
		wait for Clk_period;
		Addr <=  "0010111000110";
		Trees_din <= x"07054704";
		wait for Clk_period;
		Addr <=  "0010111000111";
		Trees_din <= x"ff811795";
		wait for Clk_period;
		Addr <=  "0010111001000";
		Trees_din <= x"00281795";
		wait for Clk_period;
		Addr <=  "0010111001001";
		Trees_din <= x"11002310";
		wait for Clk_period;
		Addr <=  "0010111001010";
		Trees_din <= x"1afcff08";
		wait for Clk_period;
		Addr <=  "0010111001011";
		Trees_din <= x"07072704";
		wait for Clk_period;
		Addr <=  "0010111001100";
		Trees_din <= x"ff751795";
		wait for Clk_period;
		Addr <=  "0010111001101";
		Trees_din <= x"00231795";
		wait for Clk_period;
		Addr <=  "0010111001110";
		Trees_din <= x"01fd2d04";
		wait for Clk_period;
		Addr <=  "0010111001111";
		Trees_din <= x"ff841795";
		wait for Clk_period;
		Addr <=  "0010111010000";
		Trees_din <= x"00531795";
		wait for Clk_period;
		Addr <=  "0010111010001";
		Trees_din <= x"0d008908";
		wait for Clk_period;
		Addr <=  "0010111010010";
		Trees_din <= x"1afc5404";
		wait for Clk_period;
		Addr <=  "0010111010011";
		Trees_din <= x"00a91795";
		wait for Clk_period;
		Addr <=  "0010111010100";
		Trees_din <= x"00081795";
		wait for Clk_period;
		Addr <=  "0010111010101";
		Trees_din <= x"15fa1c04";
		wait for Clk_period;
		Addr <=  "0010111010110";
		Trees_din <= x"ffb21795";
		wait for Clk_period;
		Addr <=  "0010111010111";
		Trees_din <= x"00511795";
		wait for Clk_period;
		Addr <=  "0010111011000";
		Trees_din <= x"0d006408";
		wait for Clk_period;
		Addr <=  "0010111011001";
		Trees_din <= x"04066204";
		wait for Clk_period;
		Addr <=  "0010111011010";
		Trees_din <= x"00fe1795";
		wait for Clk_period;
		Addr <=  "0010111011011";
		Trees_din <= x"fffa1795";
		wait for Clk_period;
		Addr <=  "0010111011100";
		Trees_din <= x"06057208";
		wait for Clk_period;
		Addr <=  "0010111011101";
		Trees_din <= x"03fb2004";
		wait for Clk_period;
		Addr <=  "0010111011110";
		Trees_din <= x"ff9d1795";
		wait for Clk_period;
		Addr <=  "0010111011111";
		Trees_din <= x"00ce1795";
		wait for Clk_period;
		Addr <=  "0010111100000";
		Trees_din <= x"0b008f04";
		wait for Clk_period;
		Addr <=  "0010111100001";
		Trees_din <= x"ff601795";
		wait for Clk_period;
		Addr <=  "0010111100010";
		Trees_din <= x"1300cc04";
		wait for Clk_period;
		Addr <=  "0010111100011";
		Trees_din <= x"fff31795";
		wait for Clk_period;
		Addr <=  "0010111100100";
		Trees_din <= x"00b71795";
		wait for Clk_period;
		Addr <=  "0010111100101";
		Trees_din <= x"11000140";
		wait for Clk_period;
		Addr <=  "0010111100110";
		Trees_din <= x"01fe5c28";
		wait for Clk_period;
		Addr <=  "0010111100111";
		Trees_din <= x"05fbb60c";
		wait for Clk_period;
		Addr <=  "0010111101000";
		Trees_din <= x"10000308";
		wait for Clk_period;
		Addr <=  "0010111101001";
		Trees_din <= x"00ff3804";
		wait for Clk_period;
		Addr <=  "0010111101010";
		Trees_din <= x"007718b9";
		wait for Clk_period;
		Addr <=  "0010111101011";
		Trees_din <= x"ffd118b9";
		wait for Clk_period;
		Addr <=  "0010111101100";
		Trees_din <= x"010618b9";
		wait for Clk_period;
		Addr <=  "0010111101101";
		Trees_din <= x"03fbe40c";
		wait for Clk_period;
		Addr <=  "0010111101110";
		Trees_din <= x"14004608";
		wait for Clk_period;
		Addr <=  "0010111101111";
		Trees_din <= x"0b00b404";
		wait for Clk_period;
		Addr <=  "0010111110000";
		Trees_din <= x"007e18b9";
		wait for Clk_period;
		Addr <=  "0010111110001";
		Trees_din <= x"ffcd18b9";
		wait for Clk_period;
		Addr <=  "0010111110010";
		Trees_din <= x"ff6318b9";
		wait for Clk_period;
		Addr <=  "0010111110011";
		Trees_din <= x"02fb3208";
		wait for Clk_period;
		Addr <=  "0010111110100";
		Trees_din <= x"02faca04";
		wait for Clk_period;
		Addr <=  "0010111110101";
		Trees_din <= x"002f18b9";
		wait for Clk_period;
		Addr <=  "0010111110110";
		Trees_din <= x"011b18b9";
		wait for Clk_period;
		Addr <=  "0010111110111";
		Trees_din <= x"02fc5b04";
		wait for Clk_period;
		Addr <=  "0010111111000";
		Trees_din <= x"ffbf18b9";
		wait for Clk_period;
		Addr <=  "0010111111001";
		Trees_din <= x"005b18b9";
		wait for Clk_period;
		Addr <=  "0010111111010";
		Trees_din <= x"0501e610";
		wait for Clk_period;
		Addr <=  "0010111111011";
		Trees_din <= x"08003f04";
		wait for Clk_period;
		Addr <=  "0010111111100";
		Trees_din <= x"004218b9";
		wait for Clk_period;
		Addr <=  "0010111111101";
		Trees_din <= x"040bc208";
		wait for Clk_period;
		Addr <=  "0010111111110";
		Trees_din <= x"0e002004";
		wait for Clk_period;
		Addr <=  "0010111111111";
		Trees_din <= x"ffe118b9";
		wait for Clk_period;
		Addr <=  "0011000000000";
		Trees_din <= x"ff7618b9";
		wait for Clk_period;
		Addr <=  "0011000000001";
		Trees_din <= x"001018b9";
		wait for Clk_period;
		Addr <=  "0011000000010";
		Trees_din <= x"07015104";
		wait for Clk_period;
		Addr <=  "0011000000011";
		Trees_din <= x"ffe418b9";
		wait for Clk_period;
		Addr <=  "0011000000100";
		Trees_din <= x"007618b9";
		wait for Clk_period;
		Addr <=  "0011000000101";
		Trees_din <= x"11000220";
		wait for Clk_period;
		Addr <=  "0011000000110";
		Trees_din <= x"1604001c";
		wait for Clk_period;
		Addr <=  "0011000000111";
		Trees_din <= x"00fd440c";
		wait for Clk_period;
		Addr <=  "0011000001000";
		Trees_din <= x"06089508";
		wait for Clk_period;
		Addr <=  "0011000001001";
		Trees_din <= x"04055c04";
		wait for Clk_period;
		Addr <=  "0011000001010";
		Trees_din <= x"00d418b9";
		wait for Clk_period;
		Addr <=  "0011000001011";
		Trees_din <= x"001818b9";
		wait for Clk_period;
		Addr <=  "0011000001100";
		Trees_din <= x"ff9118b9";
		wait for Clk_period;
		Addr <=  "0011000001101";
		Trees_din <= x"08004c08";
		wait for Clk_period;
		Addr <=  "0011000001110";
		Trees_din <= x"18006004";
		wait for Clk_period;
		Addr <=  "0011000001111";
		Trees_din <= x"ffe318b9";
		wait for Clk_period;
		Addr <=  "0011000010000";
		Trees_din <= x"ff5b18b9";
		wait for Clk_period;
		Addr <=  "0011000010001";
		Trees_din <= x"02fab104";
		wait for Clk_period;
		Addr <=  "0011000010010";
		Trees_din <= x"004d18b9";
		wait for Clk_period;
		Addr <=  "0011000010011";
		Trees_din <= x"ff9118b9";
		wait for Clk_period;
		Addr <=  "0011000010100";
		Trees_din <= x"009f18b9";
		wait for Clk_period;
		Addr <=  "0011000010101";
		Trees_din <= x"10001118";
		wait for Clk_period;
		Addr <=  "0011000010110";
		Trees_din <= x"1604000c";
		wait for Clk_period;
		Addr <=  "0011000010111";
		Trees_din <= x"05fe1f04";
		wait for Clk_period;
		Addr <=  "0011000011000";
		Trees_din <= x"ff5318b9";
		wait for Clk_period;
		Addr <=  "0011000011001";
		Trees_din <= x"03fdac04";
		wait for Clk_period;
		Addr <=  "0011000011010";
		Trees_din <= x"000918b9";
		wait for Clk_period;
		Addr <=  "0011000011011";
		Trees_din <= x"ff9518b9";
		wait for Clk_period;
		Addr <=  "0011000011100";
		Trees_din <= x"09004408";
		wait for Clk_period;
		Addr <=  "0011000011101";
		Trees_din <= x"01fed304";
		wait for Clk_period;
		Addr <=  "0011000011110";
		Trees_din <= x"ffa518b9";
		wait for Clk_period;
		Addr <=  "0011000011111";
		Trees_din <= x"00a118b9";
		wait for Clk_period;
		Addr <=  "0011000100000";
		Trees_din <= x"00c618b9";
		wait for Clk_period;
		Addr <=  "0011000100001";
		Trees_din <= x"16040010";
		wait for Clk_period;
		Addr <=  "0011000100010";
		Trees_din <= x"11000408";
		wait for Clk_period;
		Addr <=  "0011000100011";
		Trees_din <= x"00fe9104";
		wait for Clk_period;
		Addr <=  "0011000100100";
		Trees_din <= x"00cf18b9";
		wait for Clk_period;
		Addr <=  "0011000100101";
		Trees_din <= x"ffc718b9";
		wait for Clk_period;
		Addr <=  "0011000100110";
		Trees_din <= x"11000b04";
		wait for Clk_period;
		Addr <=  "0011000100111";
		Trees_din <= x"ffdb18b9";
		wait for Clk_period;
		Addr <=  "0011000101000";
		Trees_din <= x"000b18b9";
		wait for Clk_period;
		Addr <=  "0011000101001";
		Trees_din <= x"00ffa908";
		wait for Clk_period;
		Addr <=  "0011000101010";
		Trees_din <= x"05fe5404";
		wait for Clk_period;
		Addr <=  "0011000101011";
		Trees_din <= x"011818b9";
		wait for Clk_period;
		Addr <=  "0011000101100";
		Trees_din <= x"ffe518b9";
		wait for Clk_period;
		Addr <=  "0011000101101";
		Trees_din <= x"ff9018b9";
		wait for Clk_period;
		Addr <=  "0011000101110";
		Trees_din <= x"07035774";
		wait for Clk_period;
		Addr <=  "0011000101111";
		Trees_din <= x"1200503c";
		wait for Clk_period;
		Addr <=  "0011000110000";
		Trees_din <= x"1400451c";
		wait for Clk_period;
		Addr <=  "0011000110001";
		Trees_din <= x"16040010";
		wait for Clk_period;
		Addr <=  "0011000110010";
		Trees_din <= x"0e003708";
		wait for Clk_period;
		Addr <=  "0011000110011";
		Trees_din <= x"0d006704";
		wait for Clk_period;
		Addr <=  "0011000110100";
		Trees_din <= x"00721a5d";
		wait for Clk_period;
		Addr <=  "0011000110101";
		Trees_din <= x"fff61a5d";
		wait for Clk_period;
		Addr <=  "0011000110110";
		Trees_din <= x"1e027804";
		wait for Clk_period;
		Addr <=  "0011000110111";
		Trees_din <= x"ff8d1a5d";
		wait for Clk_period;
		Addr <=  "0011000111000";
		Trees_din <= x"00281a5d";
		wait for Clk_period;
		Addr <=  "0011000111001";
		Trees_din <= x"0609d108";
		wait for Clk_period;
		Addr <=  "0011000111010";
		Trees_din <= x"14004004";
		wait for Clk_period;
		Addr <=  "0011000111011";
		Trees_din <= x"00f21a5d";
		wait for Clk_period;
		Addr <=  "0011000111100";
		Trees_din <= x"002d1a5d";
		wait for Clk_period;
		Addr <=  "0011000111101";
		Trees_din <= x"ffa51a5d";
		wait for Clk_period;
		Addr <=  "0011000111110";
		Trees_din <= x"19000010";
		wait for Clk_period;
		Addr <=  "0011000111111";
		Trees_din <= x"0d006308";
		wait for Clk_period;
		Addr <=  "0011001000000";
		Trees_din <= x"0b010a04";
		wait for Clk_period;
		Addr <=  "0011001000001";
		Trees_din <= x"ffa71a5d";
		wait for Clk_period;
		Addr <=  "0011001000010";
		Trees_din <= x"007e1a5d";
		wait for Clk_period;
		Addr <=  "0011001000011";
		Trees_din <= x"1afd4304";
		wait for Clk_period;
		Addr <=  "0011001000100";
		Trees_din <= x"00c91a5d";
		wait for Clk_period;
		Addr <=  "0011001000101";
		Trees_din <= x"ffdf1a5d";
		wait for Clk_period;
		Addr <=  "0011001000110";
		Trees_din <= x"07019808";
		wait for Clk_period;
		Addr <=  "0011001000111";
		Trees_din <= x"14004504";
		wait for Clk_period;
		Addr <=  "0011001001000";
		Trees_din <= x"002e1a5d";
		wait for Clk_period;
		Addr <=  "0011001001001";
		Trees_din <= x"ff6b1a5d";
		wait for Clk_period;
		Addr <=  "0011001001010";
		Trees_din <= x"02faf804";
		wait for Clk_period;
		Addr <=  "0011001001011";
		Trees_din <= x"ff9e1a5d";
		wait for Clk_period;
		Addr <=  "0011001001100";
		Trees_din <= x"00801a5d";
		wait for Clk_period;
		Addr <=  "0011001001101";
		Trees_din <= x"00fd2018";
		wait for Clk_period;
		Addr <=  "0011001001110";
		Trees_din <= x"0d00730c";
		wait for Clk_period;
		Addr <=  "0011001001111";
		Trees_din <= x"08004f08";
		wait for Clk_period;
		Addr <=  "0011001010000";
		Trees_din <= x"0b00ce04";
		wait for Clk_period;
		Addr <=  "0011001010001";
		Trees_din <= x"ff851a5d";
		wait for Clk_period;
		Addr <=  "0011001010010";
		Trees_din <= x"00001a5d";
		wait for Clk_period;
		Addr <=  "0011001010011";
		Trees_din <= x"00501a5d";
		wait for Clk_period;
		Addr <=  "0011001010100";
		Trees_din <= x"06094508";
		wait for Clk_period;
		Addr <=  "0011001010101";
		Trees_din <= x"05fc5804";
		wait for Clk_period;
		Addr <=  "0011001010110";
		Trees_din <= x"004a1a5d";
		wait for Clk_period;
		Addr <=  "0011001010111";
		Trees_din <= x"ffce1a5d";
		wait for Clk_period;
		Addr <=  "0011001011000";
		Trees_din <= x"016a1a5d";
		wait for Clk_period;
		Addr <=  "0011001011001";
		Trees_din <= x"1b024710";
		wait for Clk_period;
		Addr <=  "0011001011010";
		Trees_din <= x"1e023d08";
		wait for Clk_period;
		Addr <=  "0011001011011";
		Trees_din <= x"1c021a04";
		wait for Clk_period;
		Addr <=  "0011001011100";
		Trees_din <= x"005b1a5d";
		wait for Clk_period;
		Addr <=  "0011001011101";
		Trees_din <= x"ff881a5d";
		wait for Clk_period;
		Addr <=  "0011001011110";
		Trees_din <= x"0b00c304";
		wait for Clk_period;
		Addr <=  "0011001011111";
		Trees_din <= x"fff01a5d";
		wait for Clk_period;
		Addr <=  "0011001100000";
		Trees_din <= x"01101a5d";
		wait for Clk_period;
		Addr <=  "0011001100001";
		Trees_din <= x"0b006308";
		wait for Clk_period;
		Addr <=  "0011001100010";
		Trees_din <= x"19000104";
		wait for Clk_period;
		Addr <=  "0011001100011";
		Trees_din <= x"ffce1a5d";
		wait for Clk_period;
		Addr <=  "0011001100100";
		Trees_din <= x"00c01a5d";
		wait for Clk_period;
		Addr <=  "0011001100101";
		Trees_din <= x"10019204";
		wait for Clk_period;
		Addr <=  "0011001100110";
		Trees_din <= x"ff651a5d";
		wait for Clk_period;
		Addr <=  "0011001100111";
		Trees_din <= x"ffec1a5d";
		wait for Clk_period;
		Addr <=  "0011001101000";
		Trees_din <= x"1e025020";
		wait for Clk_period;
		Addr <=  "0011001101001";
		Trees_din <= x"1d024410";
		wait for Clk_period;
		Addr <=  "0011001101010";
		Trees_din <= x"01fdb608";
		wait for Clk_period;
		Addr <=  "0011001101011";
		Trees_din <= x"03fc0b04";
		wait for Clk_period;
		Addr <=  "0011001101100";
		Trees_din <= x"ff781a5d";
		wait for Clk_period;
		Addr <=  "0011001101101";
		Trees_din <= x"00111a5d";
		wait for Clk_period;
		Addr <=  "0011001101110";
		Trees_din <= x"0408c104";
		wait for Clk_period;
		Addr <=  "0011001101111";
		Trees_din <= x"00961a5d";
		wait for Clk_period;
		Addr <=  "0011001110000";
		Trees_din <= x"ffb81a5d";
		wait for Clk_period;
		Addr <=  "0011001110001";
		Trees_din <= x"06008e08";
		wait for Clk_period;
		Addr <=  "0011001110010";
		Trees_din <= x"05fd4204";
		wait for Clk_period;
		Addr <=  "0011001110011";
		Trees_din <= x"ffd41a5d";
		wait for Clk_period;
		Addr <=  "0011001110100";
		Trees_din <= x"00751a5d";
		wait for Clk_period;
		Addr <=  "0011001110101";
		Trees_din <= x"17040004";
		wait for Clk_period;
		Addr <=  "0011001110110";
		Trees_din <= x"00d31a5d";
		wait for Clk_period;
		Addr <=  "0011001110111";
		Trees_din <= x"003c1a5d";
		wait for Clk_period;
		Addr <=  "0011001111000";
		Trees_din <= x"19000120";
		wait for Clk_period;
		Addr <=  "0011001111001";
		Trees_din <= x"0c003a10";
		wait for Clk_period;
		Addr <=  "0011001111010";
		Trees_din <= x"0c000a08";
		wait for Clk_period;
		Addr <=  "0011001111011";
		Trees_din <= x"14004604";
		wait for Clk_period;
		Addr <=  "0011001111100";
		Trees_din <= x"009b1a5d";
		wait for Clk_period;
		Addr <=  "0011001111101";
		Trees_din <= x"ffa81a5d";
		wait for Clk_period;
		Addr <=  "0011001111110";
		Trees_din <= x"00ff3804";
		wait for Clk_period;
		Addr <=  "0011001111111";
		Trees_din <= x"fff91a5d";
		wait for Clk_period;
		Addr <=  "0011010000000";
		Trees_din <= x"ff5f1a5d";
		wait for Clk_period;
		Addr <=  "0011010000001";
		Trees_din <= x"0f008908";
		wait for Clk_period;
		Addr <=  "0011010000010";
		Trees_din <= x"09003b04";
		wait for Clk_period;
		Addr <=  "0011010000011";
		Trees_din <= x"00991a5d";
		wait for Clk_period;
		Addr <=  "0011010000100";
		Trees_din <= x"00261a5d";
		wait for Clk_period;
		Addr <=  "0011010000101";
		Trees_din <= x"05fd8904";
		wait for Clk_period;
		Addr <=  "0011010000110";
		Trees_din <= x"ff7c1a5d";
		wait for Clk_period;
		Addr <=  "0011010000111";
		Trees_din <= x"00231a5d";
		wait for Clk_period;
		Addr <=  "0011010001000";
		Trees_din <= x"07054710";
		wait for Clk_period;
		Addr <=  "0011010001001";
		Trees_din <= x"18004c08";
		wait for Clk_period;
		Addr <=  "0011010001010";
		Trees_din <= x"04057c04";
		wait for Clk_period;
		Addr <=  "0011010001011";
		Trees_din <= x"007b1a5d";
		wait for Clk_period;
		Addr <=  "0011010001100";
		Trees_din <= x"fff61a5d";
		wait for Clk_period;
		Addr <=  "0011010001101";
		Trees_din <= x"1703e004";
		wait for Clk_period;
		Addr <=  "0011010001110";
		Trees_din <= x"ff671a5d";
		wait for Clk_period;
		Addr <=  "0011010001111";
		Trees_din <= x"00081a5d";
		wait for Clk_period;
		Addr <=  "0011010010000";
		Trees_din <= x"03fc7808";
		wait for Clk_period;
		Addr <=  "0011010010001";
		Trees_din <= x"00ffd204";
		wait for Clk_period;
		Addr <=  "0011010010010";
		Trees_din <= x"005f1a5d";
		wait for Clk_period;
		Addr <=  "0011010010011";
		Trees_din <= x"ffb21a5d";
		wait for Clk_period;
		Addr <=  "0011010010100";
		Trees_din <= x"00036a04";
		wait for Clk_period;
		Addr <=  "0011010010101";
		Trees_din <= x"00921a5d";
		wait for Clk_period;
		Addr <=  "0011010010110";
		Trees_din <= x"001a1a5d";
		wait for Clk_period;
		Addr <=  "0011010010111";
		Trees_din <= x"07072754";
		wait for Clk_period;
		Addr <=  "0011010011000";
		Trees_din <= x"0e001f28";
		wait for Clk_period;
		Addr <=  "0011010011001";
		Trees_din <= x"0f009b20";
		wait for Clk_period;
		Addr <=  "0011010011010";
		Trees_din <= x"00fe7e10";
		wait for Clk_period;
		Addr <=  "0011010011011";
		Trees_din <= x"00fdc408";
		wait for Clk_period;
		Addr <=  "0011010011100";
		Trees_din <= x"0603f604";
		wait for Clk_period;
		Addr <=  "0011010011101";
		Trees_din <= x"00631b59";
		wait for Clk_period;
		Addr <=  "0011010011110";
		Trees_din <= x"ffc71b59";
		wait for Clk_period;
		Addr <=  "0011010011111";
		Trees_din <= x"05fdb604";
		wait for Clk_period;
		Addr <=  "0011010100000";
		Trees_din <= x"003c1b59";
		wait for Clk_period;
		Addr <=  "0011010100001";
		Trees_din <= x"00e31b59";
		wait for Clk_period;
		Addr <=  "0011010100010";
		Trees_din <= x"0a00aa08";
		wait for Clk_period;
		Addr <=  "0011010100011";
		Trees_din <= x"16040004";
		wait for Clk_period;
		Addr <=  "0011010100100";
		Trees_din <= x"ffbd1b59";
		wait for Clk_period;
		Addr <=  "0011010100101";
		Trees_din <= x"007b1b59";
		wait for Clk_period;
		Addr <=  "0011010100110";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "0011010100111";
		Trees_din <= x"ffb61b59";
		wait for Clk_period;
		Addr <=  "0011010101000";
		Trees_din <= x"00981b59";
		wait for Clk_period;
		Addr <=  "0011010101001";
		Trees_din <= x"0601e804";
		wait for Clk_period;
		Addr <=  "0011010101010";
		Trees_din <= x"00151b59";
		wait for Clk_period;
		Addr <=  "0011010101011";
		Trees_din <= x"ff7b1b59";
		wait for Clk_period;
		Addr <=  "0011010101100";
		Trees_din <= x"040a1520";
		wait for Clk_period;
		Addr <=  "0011010101101";
		Trees_din <= x"00fd4410";
		wait for Clk_period;
		Addr <=  "0011010101110";
		Trees_din <= x"14003608";
		wait for Clk_period;
		Addr <=  "0011010101111";
		Trees_din <= x"02fb2804";
		wait for Clk_period;
		Addr <=  "0011010110000";
		Trees_din <= x"ff681b59";
		wait for Clk_period;
		Addr <=  "0011010110001";
		Trees_din <= x"00391b59";
		wait for Clk_period;
		Addr <=  "0011010110010";
		Trees_din <= x"0f006a04";
		wait for Clk_period;
		Addr <=  "0011010110011";
		Trees_din <= x"ffc31b59";
		wait for Clk_period;
		Addr <=  "0011010110100";
		Trees_din <= x"004d1b59";
		wait for Clk_period;
		Addr <=  "0011010110101";
		Trees_din <= x"03fcf208";
		wait for Clk_period;
		Addr <=  "0011010110110";
		Trees_din <= x"0001c404";
		wait for Clk_period;
		Addr <=  "0011010110111";
		Trees_din <= x"00101b59";
		wait for Clk_period;
		Addr <=  "0011010111000";
		Trees_din <= x"ff921b59";
		wait for Clk_period;
		Addr <=  "0011010111001";
		Trees_din <= x"03fdac04";
		wait for Clk_period;
		Addr <=  "0011010111010";
		Trees_din <= x"ffa91b59";
		wait for Clk_period;
		Addr <=  "0011010111011";
		Trees_din <= x"fffb1b59";
		wait for Clk_period;
		Addr <=  "0011010111100";
		Trees_din <= x"10030a08";
		wait for Clk_period;
		Addr <=  "0011010111101";
		Trees_din <= x"02fdb404";
		wait for Clk_period;
		Addr <=  "0011010111110";
		Trees_din <= x"ff721b59";
		wait for Clk_period;
		Addr <=  "0011010111111";
		Trees_din <= x"00081b59";
		wait for Clk_period;
		Addr <=  "0011011000000";
		Trees_din <= x"00321b59";
		wait for Clk_period;
		Addr <=  "0011011000001";
		Trees_din <= x"02f8fa10";
		wait for Clk_period;
		Addr <=  "0011011000010";
		Trees_din <= x"17037c08";
		wait for Clk_period;
		Addr <=  "0011011000011";
		Trees_din <= x"01fdbf04";
		wait for Clk_period;
		Addr <=  "0011011000100";
		Trees_din <= x"005d1b59";
		wait for Clk_period;
		Addr <=  "0011011000101";
		Trees_din <= x"fff01b59";
		wait for Clk_period;
		Addr <=  "0011011000110";
		Trees_din <= x"05fcf004";
		wait for Clk_period;
		Addr <=  "0011011000111";
		Trees_din <= x"ff701b59";
		wait for Clk_period;
		Addr <=  "0011011001000";
		Trees_din <= x"000e1b59";
		wait for Clk_period;
		Addr <=  "0011011001001";
		Trees_din <= x"0100ff14";
		wait for Clk_period;
		Addr <=  "0011011001010";
		Trees_din <= x"05fbbf0c";
		wait for Clk_period;
		Addr <=  "0011011001011";
		Trees_din <= x"0b00b304";
		wait for Clk_period;
		Addr <=  "0011011001100";
		Trees_din <= x"00721b59";
		wait for Clk_period;
		Addr <=  "0011011001101";
		Trees_din <= x"02faf204";
		wait for Clk_period;
		Addr <=  "0011011001110";
		Trees_din <= x"ffa81b59";
		wait for Clk_period;
		Addr <=  "0011011001111";
		Trees_din <= x"00281b59";
		wait for Clk_period;
		Addr <=  "0011011010000";
		Trees_din <= x"13008804";
		wait for Clk_period;
		Addr <=  "0011011010001";
		Trees_din <= x"001f1b59";
		wait for Clk_period;
		Addr <=  "0011011010010";
		Trees_din <= x"008d1b59";
		wait for Clk_period;
		Addr <=  "0011011010011";
		Trees_din <= x"02fd4d04";
		wait for Clk_period;
		Addr <=  "0011011010100";
		Trees_din <= x"ffa81b59";
		wait for Clk_period;
		Addr <=  "0011011010101";
		Trees_din <= x"005f1b59";
		wait for Clk_period;
		Addr <=  "0011011010110";
		Trees_din <= x"0703572c";
		wait for Clk_period;
		Addr <=  "0011011010111";
		Trees_din <= x"02f91404";
		wait for Clk_period;
		Addr <=  "0011011011000";
		Trees_din <= x"ff731c4d";
		wait for Clk_period;
		Addr <=  "0011011011001";
		Trees_din <= x"0409321c";
		wait for Clk_period;
		Addr <=  "0011011011010";
		Trees_din <= x"0408ab10";
		wait for Clk_period;
		Addr <=  "0011011011011";
		Trees_din <= x"12005008";
		wait for Clk_period;
		Addr <=  "0011011011100";
		Trees_din <= x"0e004404";
		wait for Clk_period;
		Addr <=  "0011011011101";
		Trees_din <= x"00011c4d";
		wait for Clk_period;
		Addr <=  "0011011011110";
		Trees_din <= x"00611c4d";
		wait for Clk_period;
		Addr <=  "0011011011111";
		Trees_din <= x"00fd2004";
		wait for Clk_period;
		Addr <=  "0011011100000";
		Trees_din <= x"00581c4d";
		wait for Clk_period;
		Addr <=  "0011011100001";
		Trees_din <= x"ffc51c4d";
		wait for Clk_period;
		Addr <=  "0011011100010";
		Trees_din <= x"05fce508";
		wait for Clk_period;
		Addr <=  "0011011100011";
		Trees_din <= x"0c01db04";
		wait for Clk_period;
		Addr <=  "0011011100100";
		Trees_din <= x"010c1c4d";
		wait for Clk_period;
		Addr <=  "0011011100101";
		Trees_din <= x"ffd71c4d";
		wait for Clk_period;
		Addr <=  "0011011100110";
		Trees_din <= x"ff871c4d";
		wait for Clk_period;
		Addr <=  "0011011100111";
		Trees_din <= x"07028104";
		wait for Clk_period;
		Addr <=  "0011011101000";
		Trees_din <= x"ff761c4d";
		wait for Clk_period;
		Addr <=  "0011011101001";
		Trees_din <= x"1603f504";
		wait for Clk_period;
		Addr <=  "0011011101010";
		Trees_din <= x"003e1c4d";
		wait for Clk_period;
		Addr <=  "0011011101011";
		Trees_din <= x"00041c4d";
		wait for Clk_period;
		Addr <=  "0011011101100";
		Trees_din <= x"1e02501c";
		wait for Clk_period;
		Addr <=  "0011011101101";
		Trees_din <= x"1d024410";
		wait for Clk_period;
		Addr <=  "0011011101110";
		Trees_din <= x"01fdb608";
		wait for Clk_period;
		Addr <=  "0011011101111";
		Trees_din <= x"0705d204";
		wait for Clk_period;
		Addr <=  "0011011110000";
		Trees_din <= x"ff791c4d";
		wait for Clk_period;
		Addr <=  "0011011110001";
		Trees_din <= x"000d1c4d";
		wait for Clk_period;
		Addr <=  "0011011110010";
		Trees_din <= x"01ffcd04";
		wait for Clk_period;
		Addr <=  "0011011110011";
		Trees_din <= x"008e1c4d";
		wait for Clk_period;
		Addr <=  "0011011110100";
		Trees_din <= x"ffca1c4d";
		wait for Clk_period;
		Addr <=  "0011011110101";
		Trees_din <= x"18008b08";
		wait for Clk_period;
		Addr <=  "0011011110110";
		Trees_din <= x"06fe9d04";
		wait for Clk_period;
		Addr <=  "0011011110111";
		Trees_din <= x"003e1c4d";
		wait for Clk_period;
		Addr <=  "0011011111000";
		Trees_din <= x"00b81c4d";
		wait for Clk_period;
		Addr <=  "0011011111001";
		Trees_din <= x"00201c4d";
		wait for Clk_period;
		Addr <=  "0011011111010";
		Trees_din <= x"18005314";
		wait for Clk_period;
		Addr <=  "0011011111011";
		Trees_din <= x"0d00ab0c";
		wait for Clk_period;
		Addr <=  "0011011111100";
		Trees_din <= x"06fdfe08";
		wait for Clk_period;
		Addr <=  "0011011111101";
		Trees_din <= x"15f7c104";
		wait for Clk_period;
		Addr <=  "0011011111110";
		Trees_din <= x"ffa51c4d";
		wait for Clk_period;
		Addr <=  "0011011111111";
		Trees_din <= x"004b1c4d";
		wait for Clk_period;
		Addr <=  "0011100000000";
		Trees_din <= x"00b41c4d";
		wait for Clk_period;
		Addr <=  "0011100000001";
		Trees_din <= x"02fa1604";
		wait for Clk_period;
		Addr <=  "0011100000010";
		Trees_din <= x"ff881c4d";
		wait for Clk_period;
		Addr <=  "0011100000011";
		Trees_din <= x"fff71c4d";
		wait for Clk_period;
		Addr <=  "0011100000100";
		Trees_din <= x"19000110";
		wait for Clk_period;
		Addr <=  "0011100000101";
		Trees_din <= x"0c003a08";
		wait for Clk_period;
		Addr <=  "0011100000110";
		Trees_din <= x"0c000e04";
		wait for Clk_period;
		Addr <=  "0011100000111";
		Trees_din <= x"001a1c4d";
		wait for Clk_period;
		Addr <=  "0011100001000";
		Trees_din <= x"ff831c4d";
		wait for Clk_period;
		Addr <=  "0011100001001";
		Trees_din <= x"1300c004";
		wait for Clk_period;
		Addr <=  "0011100001010";
		Trees_din <= x"00371c4d";
		wait for Clk_period;
		Addr <=  "0011100001011";
		Trees_din <= x"ffb91c4d";
		wait for Clk_period;
		Addr <=  "0011100001100";
		Trees_din <= x"07054708";
		wait for Clk_period;
		Addr <=  "0011100001101";
		Trees_din <= x"04044104";
		wait for Clk_period;
		Addr <=  "0011100001110";
		Trees_din <= x"00001c4d";
		wait for Clk_period;
		Addr <=  "0011100001111";
		Trees_din <= x"ff681c4d";
		wait for Clk_period;
		Addr <=  "0011100010000";
		Trees_din <= x"1e027804";
		wait for Clk_period;
		Addr <=  "0011100010001";
		Trees_din <= x"00511c4d";
		wait for Clk_period;
		Addr <=  "0011100010010";
		Trees_din <= x"ffd21c4d";
		wait for Clk_period;
		Addr <=  "0011100010011";
		Trees_din <= x"15f6ca0c";
		wait for Clk_period;
		Addr <=  "0011100010100";
		Trees_din <= x"1e020904";
		wait for Clk_period;
		Addr <=  "0011100010101";
		Trees_din <= x"003d1d09";
		wait for Clk_period;
		Addr <=  "0011100010110";
		Trees_din <= x"08004d04";
		wait for Clk_period;
		Addr <=  "0011100010111";
		Trees_din <= x"ff6f1d09";
		wait for Clk_period;
		Addr <=  "0011100011000";
		Trees_din <= x"ffff1d09";
		wait for Clk_period;
		Addr <=  "0011100011001";
		Trees_din <= x"15f6fc20";
		wait for Clk_period;
		Addr <=  "0011100011010";
		Trees_din <= x"06099918";
		wait for Clk_period;
		Addr <=  "0011100011011";
		Trees_din <= x"06077b10";
		wait for Clk_period;
		Addr <=  "0011100011100";
		Trees_din <= x"01fd9608";
		wait for Clk_period;
		Addr <=  "0011100011101";
		Trees_din <= x"0a000904";
		wait for Clk_period;
		Addr <=  "0011100011110";
		Trees_din <= x"ffe11d09";
		wait for Clk_period;
		Addr <=  "0011100011111";
		Trees_din <= x"ff8c1d09";
		wait for Clk_period;
		Addr <=  "0011100100000";
		Trees_din <= x"03fd1304";
		wait for Clk_period;
		Addr <=  "0011100100001";
		Trees_din <= x"fff11d09";
		wait for Clk_period;
		Addr <=  "0011100100010";
		Trees_din <= x"00811d09";
		wait for Clk_period;
		Addr <=  "0011100100011";
		Trees_din <= x"0b00d204";
		wait for Clk_period;
		Addr <=  "0011100100100";
		Trees_din <= x"00191d09";
		wait for Clk_period;
		Addr <=  "0011100100101";
		Trees_din <= x"01341d09";
		wait for Clk_period;
		Addr <=  "0011100100110";
		Trees_din <= x"0d005104";
		wait for Clk_period;
		Addr <=  "0011100100111";
		Trees_din <= x"00281d09";
		wait for Clk_period;
		Addr <=  "0011100101000";
		Trees_din <= x"ff8e1d09";
		wait for Clk_period;
		Addr <=  "0011100101001";
		Trees_din <= x"07015b14";
		wait for Clk_period;
		Addr <=  "0011100101010";
		Trees_din <= x"1300f810";
		wait for Clk_period;
		Addr <=  "0011100101011";
		Trees_din <= x"0f008808";
		wait for Clk_period;
		Addr <=  "0011100101100";
		Trees_din <= x"09003f04";
		wait for Clk_period;
		Addr <=  "0011100101101";
		Trees_din <= x"ffd01d09";
		wait for Clk_period;
		Addr <=  "0011100101110";
		Trees_din <= x"00071d09";
		wait for Clk_period;
		Addr <=  "0011100101111";
		Trees_din <= x"09003d04";
		wait for Clk_period;
		Addr <=  "0011100110000";
		Trees_din <= x"00921d09";
		wait for Clk_period;
		Addr <=  "0011100110001";
		Trees_din <= x"fff61d09";
		wait for Clk_period;
		Addr <=  "0011100110010";
		Trees_din <= x"ff781d09";
		wait for Clk_period;
		Addr <=  "0011100110011";
		Trees_din <= x"02face10";
		wait for Clk_period;
		Addr <=  "0011100110100";
		Trees_din <= x"03fc2208";
		wait for Clk_period;
		Addr <=  "0011100110101";
		Trees_din <= x"02fa2e04";
		wait for Clk_period;
		Addr <=  "0011100110110";
		Trees_din <= x"002f1d09";
		wait for Clk_period;
		Addr <=  "0011100110111";
		Trees_din <= x"ffd71d09";
		wait for Clk_period;
		Addr <=  "0011100111000";
		Trees_din <= x"04041504";
		wait for Clk_period;
		Addr <=  "0011100111001";
		Trees_din <= x"00251d09";
		wait for Clk_period;
		Addr <=  "0011100111010";
		Trees_din <= x"ffb81d09";
		wait for Clk_period;
		Addr <=  "0011100111011";
		Trees_din <= x"0f008508";
		wait for Clk_period;
		Addr <=  "0011100111100";
		Trees_din <= x"08003f04";
		wait for Clk_period;
		Addr <=  "0011100111101";
		Trees_din <= x"ffd71d09";
		wait for Clk_period;
		Addr <=  "0011100111110";
		Trees_din <= x"00451d09";
		wait for Clk_period;
		Addr <=  "0011100111111";
		Trees_din <= x"0605c304";
		wait for Clk_period;
		Addr <=  "0011101000000";
		Trees_din <= x"00141d09";
		wait for Clk_period;
		Addr <=  "0011101000001";
		Trees_din <= x"ff801d09";
		wait for Clk_period;
		Addr <=  "0011101000010";
		Trees_din <= x"0000001f";
		wait for Clk_period;

        -- Reset valid flag
        Valid_node <= '0';
        wait for Clk_period; 
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111100011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101010110";
        wait for Clk_period; 
        Features_din <= "1111111001110111";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000000110000010";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "1111111000111000";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000001000111010";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000100110010";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000011001010";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111100001111000";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000000011001011";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111101100010100";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111001010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111001111011";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000000111010100";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "1111111001000000";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000001001010010";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000100001111";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "0000000110101100";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000011000110";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111100000001111";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001100010101";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101110101011";
        wait for Clk_period; 
        Features_din <= "0000001001110101";
        wait for Clk_period; 
        Features_din <= "0000001001110101";
        wait for Clk_period; 
        Features_din <= "0000001001110101";
        wait for Clk_period; 
        Features_din <= "0000001001110101";
        wait for Clk_period; 
        Features_din <= "0000001001110101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110110100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111001010000";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "0000000110010000";
        wait for Clk_period; 
        Features_din <= "0000000011011010";
        wait for Clk_period; 
        Features_din <= "1111111001001100";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000000011010101";
        wait for Clk_period; 
        Features_din <= "0000000011100000";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000000100000110";
        wait for Clk_period; 
        Features_din <= "0000000100010110";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000011110010";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111101000111000";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "1111100100101010";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(6, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111010000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111000110101";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "0000000110011111";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "1111111000101101";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000010101100";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111011101001110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110011111110";
        wait for Clk_period; 
        Features_din <= "0000001001010111";
        wait for Clk_period; 
        Features_din <= "0000001001010111";
        wait for Clk_period; 
        Features_din <= "0000001001010111";
        wait for Clk_period; 
        Features_din <= "0000001001010111";
        wait for Clk_period; 
        Features_din <= "0000001001010111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(5, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111010010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111001101011";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000000110000110";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "1111111001101110";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "0000000011111000";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111011101110010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111110010110110";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111001010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111000111011";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "0000000110000011";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "1111111001101001";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000011011111";
        wait for Clk_period; 
        Features_din <= "0000001011111100";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000001000101010";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111100001001010";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001010011010";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101101010011";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111010001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100110000";
        wait for Clk_period; 
        Features_din <= "1111111001011011";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "0000000010101101";
        wait for Clk_period; 
        Features_din <= "0000000101100101";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "1111111001000100";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000011011111";
        wait for Clk_period; 
        Features_din <= "0000000110000110";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000011000101";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111011110011000";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110001101111";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(5, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111000111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111001010101";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "0000000110111010";
        wait for Clk_period; 
        Features_din <= "0000000010111000";
        wait for Clk_period; 
        Features_din <= "1111111001001100";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "1111011111101111";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101111011101";
        wait for Clk_period; 
        Features_din <= "0000001001110001";
        wait for Clk_period; 
        Features_din <= "0000001001110001";
        wait for Clk_period; 
        Features_din <= "0000001001110001";
        wait for Clk_period; 
        Features_din <= "0000001001110001";
        wait for Clk_period; 
        Features_din <= "0000001001110001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111100000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111001101000";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000101110011";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "1111111000110111";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000111000100";
        wait for Clk_period; 
        Features_din <= "0000000011111011";
        wait for Clk_period; 
        Features_din <= "0000001001001000";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000011110001";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111100001000111";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001011000101";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111101101011000";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110101110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111111001100001";
        wait for Clk_period; 
        Features_din <= "1111111111101011";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000110011000";
        wait for Clk_period; 
        Features_din <= "0000000011011010";
        wait for Clk_period; 
        Features_din <= "1111111000110101";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111011100110100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110100110101";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111101010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111001100000";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000000110111011";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "1111111001011110";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000011011011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000000011001110";
        wait for Clk_period; 
        Features_din <= "0000001011111010";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000110011010";
        wait for Clk_period; 
        Features_din <= "0000001010001010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "1111100111110001";
        wait for Clk_period; 
        Features_din <= "0000010011011000";
        wait for Clk_period; 
        Features_din <= "1111110110010111";
        wait for Clk_period; 
        Features_din <= "0000010111011101";
        wait for Clk_period; 
        Features_din <= "1111110100101010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111000110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111001101111";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "0000000101100110";
        wait for Clk_period; 
        Features_din <= "0000000010111101";
        wait for Clk_period; 
        Features_din <= "1111111000110110";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000000100000000";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111011100000111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110110011110";
        wait for Clk_period; 
        Features_din <= "0000001001000101";
        wait for Clk_period; 
        Features_din <= "0000001001000101";
        wait for Clk_period; 
        Features_din <= "0000001001000101";
        wait for Clk_period; 
        Features_din <= "0000001001000101";
        wait for Clk_period; 
        Features_din <= "0000001001000101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111010101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "1111111001001011";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "0000000110011010";
        wait for Clk_period; 
        Features_din <= "0000000011100111";
        wait for Clk_period; 
        Features_din <= "1111111001001011";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000011010101";
        wait for Clk_period; 
        Features_din <= "0000000010110010";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111011101011000";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110011101010";
        wait for Clk_period; 
        Features_din <= "0000001001011001";
        wait for Clk_period; 
        Features_din <= "0000001001011001";
        wait for Clk_period; 
        Features_din <= "0000001001011001";
        wait for Clk_period; 
        Features_din <= "0000001001011001";
        wait for Clk_period; 
        Features_din <= "0000001001011001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111001000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100110010";
        wait for Clk_period; 
        Features_din <= "1111111000111000";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "0000000110001100";
        wait for Clk_period; 
        Features_din <= "0000000100001010";
        wait for Clk_period; 
        Features_din <= "1111111001101101";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000000011101100";
        wait for Clk_period; 
        Features_din <= "0000000100000111";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "1111011110010010";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111110001111100";
        wait for Clk_period; 
        Features_din <= "0000001001100100";
        wait for Clk_period; 
        Features_din <= "0000001001100100";
        wait for Clk_period; 
        Features_din <= "0000001001100100";
        wait for Clk_period; 
        Features_din <= "0000001001100100";
        wait for Clk_period; 
        Features_din <= "0000001001100100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110110110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101001111";
        wait for Clk_period; 
        Features_din <= "1111111000110111";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "0000000011001101";
        wait for Clk_period; 
        Features_din <= "0000000101111000";
        wait for Clk_period; 
        Features_din <= "0000000011110000";
        wait for Clk_period; 
        Features_din <= "1111111001100100";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000000011011111";
        wait for Clk_period; 
        Features_din <= "0000000011101010";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111011011101100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110111100001";
        wait for Clk_period; 
        Features_din <= "0000001000111101";
        wait for Clk_period; 
        Features_din <= "0000001000111101";
        wait for Clk_period; 
        Features_din <= "0000001000111101";
        wait for Clk_period; 
        Features_din <= "0000001000111101";
        wait for Clk_period; 
        Features_din <= "0000001000111101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110111111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111000111110";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "0000000110011011";
        wait for Clk_period; 
        Features_din <= "0000000011001001";
        wait for Clk_period; 
        Features_din <= "1111111000110101";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000001000101010";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "0000000011111010";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111011101000010";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001001010010";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110100011001";
        wait for Clk_period; 
        Features_din <= "0000001001010100";
        wait for Clk_period; 
        Features_din <= "0000001001010100";
        wait for Clk_period; 
        Features_din <= "0000001001010100";
        wait for Clk_period; 
        Features_din <= "0000001001010100";
        wait for Clk_period; 
        Features_din <= "0000001001010100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111000111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111000101001";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000110010010";
        wait for Clk_period; 
        Features_din <= "0000000011100011";
        wait for Clk_period; 
        Features_din <= "1111111001011001";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000100001011";
        wait for Clk_period; 
        Features_din <= "0000000011100010";
        wait for Clk_period; 
        Features_din <= "0000000011110011";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000000011001100";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000010111100";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111011111010111";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110000000011";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111011100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101010011";
        wait for Clk_period; 
        Features_din <= "1111111000101111";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "0000000101101110";
        wait for Clk_period; 
        Features_din <= "0000000011100101";
        wait for Clk_period; 
        Features_din <= "1111111001100000";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000011101100";
        wait for Clk_period; 
        Features_din <= "0000000110011110";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "0000000011100111";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111100000101110";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111101101111011";
        wait for Clk_period; 
        Features_din <= "0000001001111000";
        wait for Clk_period; 
        Features_din <= "0000001001111000";
        wait for Clk_period; 
        Features_din <= "0000001001111000";
        wait for Clk_period; 
        Features_din <= "0000001001111000";
        wait for Clk_period; 
        Features_din <= "0000001001111000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110110101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111001100000";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000000110000111";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "1111111001111011";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "0000000100000011";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111011110000010";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110010011000";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111110001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "1111111000111101";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "0000000101011011";
        wait for Clk_period; 
        Features_din <= "0000000011100000";
        wait for Clk_period; 
        Features_din <= "1111111001011100";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000011100101";
        wait for Clk_period; 
        Features_din <= "0000000011101110";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111011110011000";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110001101111";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111000000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111000100010";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "0000000101011011";
        wait for Clk_period; 
        Features_din <= "0000000011011101";
        wait for Clk_period; 
        Features_din <= "1111111001111101";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000011110010";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "1111011101001110";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111110011111111";
        wait for Clk_period; 
        Features_din <= "0000001001010111";
        wait for Clk_period; 
        Features_din <= "0000001001010111";
        wait for Clk_period; 
        Features_din <= "0000001001010111";
        wait for Clk_period; 
        Features_din <= "0000001001010111";
        wait for Clk_period; 
        Features_din <= "0000001001010111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110110101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111001001011";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "0000000110010010";
        wait for Clk_period; 
        Features_din <= "0000000011010011";
        wait for Clk_period; 
        Features_din <= "1111111001000100";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000110100000";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "0000001001010011";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111011100111110";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001011010010";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110100100010";
        wait for Clk_period; 
        Features_din <= "0000001001010011";
        wait for Clk_period; 
        Features_din <= "0000001001010011";
        wait for Clk_period; 
        Features_din <= "0000001001010011";
        wait for Clk_period; 
        Features_din <= "0000001001010011";
        wait for Clk_period; 
        Features_din <= "0000001001010011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111110101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111001000101";
        wait for Clk_period; 
        Features_din <= "1111111111100010";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000101110001";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "1111111001011111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "0000000011100001";
        wait for Clk_period; 
        Features_din <= "0000000101101110";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000011001110";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111100001101011";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111101100100101";
        wait for Clk_period; 
        Features_din <= "0000001001111101";
        wait for Clk_period; 
        Features_din <= "0000001001111101";
        wait for Clk_period; 
        Features_din <= "0000001001111101";
        wait for Clk_period; 
        Features_din <= "0000001001111101";
        wait for Clk_period; 
        Features_din <= "0000001001111101";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111010101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111001111101";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000110010111";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "1111111000101000";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000011100111";
        wait for Clk_period; 
        Features_din <= "0000000101010111";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000011000000";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111011110100001";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110001100000";
        wait for Clk_period; 
        Features_din <= "0000001001100110";
        wait for Clk_period; 
        Features_din <= "0000001001100110";
        wait for Clk_period; 
        Features_din <= "0000001001100110";
        wait for Clk_period; 
        Features_din <= "0000001001100110";
        wait for Clk_period; 
        Features_din <= "0000001001100110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(6, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110111110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111001101100";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000110101000";
        wait for Clk_period; 
        Features_din <= "0000000011001100";
        wait for Clk_period; 
        Features_din <= "1111111001010110";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000011111100";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111100001001000";
        wait for Clk_period; 
        Features_din <= "0000000011101100";
        wait for Clk_period; 
        Features_din <= "0000000011100011";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101101010110";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111011001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111001011000";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "0000000110000101";
        wait for Clk_period; 
        Features_din <= "0000000011100001";
        wait for Clk_period; 
        Features_din <= "1111111001011001";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000000011100001";
        wait for Clk_period; 
        Features_din <= "0000000101101001";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111100011000000";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111101010110101";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111010100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111001000001";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "0000000011000100";
        wait for Clk_period; 
        Features_din <= "0000000101110011";
        wait for Clk_period; 
        Features_din <= "0000000011100111";
        wait for Clk_period; 
        Features_din <= "1111111001001011";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000011100100";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010111100";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111011111001101";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111110000010101";
        wait for Clk_period; 
        Features_din <= "0000001001101101";
        wait for Clk_period; 
        Features_din <= "0000001001101101";
        wait for Clk_period; 
        Features_din <= "0000001001101101";
        wait for Clk_period; 
        Features_din <= "0000001001101101";
        wait for Clk_period; 
        Features_din <= "0000001001101101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111011001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101011111";
        wait for Clk_period; 
        Features_din <= "1111111001111000";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "0000000101110100";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "1111111001001111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000011101010";
        wait for Clk_period; 
        Features_din <= "0000000011011110";
        wait for Clk_period; 
        Features_din <= "0000000011011101";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000011000110";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111011110001000";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110010001110";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111001011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111001011100";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "0000000101110011";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "1111111001001110";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "0000000110111110";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000000101011111";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000011001000";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111100010111110";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111101010111001";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110111011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111001010100";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "0000000011001111";
        wait for Clk_period; 
        Features_din <= "0000000110000011";
        wait for Clk_period; 
        Features_din <= "0000000100000011";
        wait for Clk_period; 
        Features_din <= "1111111001110010";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "0000000011101000";
        wait for Clk_period; 
        Features_din <= "0000000100111001";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111011110111001";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111110000110110";
        wait for Clk_period; 
        Features_din <= "0000001001101010";
        wait for Clk_period; 
        Features_din <= "0000001001101010";
        wait for Clk_period; 
        Features_din <= "0000001001101010";
        wait for Clk_period; 
        Features_din <= "0000001001101010";
        wait for Clk_period; 
        Features_din <= "0000001001101010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111100111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111001011111";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000110110000";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "1111111000100101";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000010111100";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111011110101100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111110001001100";
        wait for Clk_period; 
        Features_din <= "0000001001101000";
        wait for Clk_period; 
        Features_din <= "0000001001101000";
        wait for Clk_period; 
        Features_din <= "0000001001101000";
        wait for Clk_period; 
        Features_din <= "0000001001101000";
        wait for Clk_period; 
        Features_din <= "0000001001101000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110111110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111001000010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "0000000110011000";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "1111111001000100";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000100011101";
        wait for Clk_period; 
        Features_din <= "0000000101110101";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000010111101";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111100000110011";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111101101110100";
        wait for Clk_period; 
        Features_din <= "0000001001111000";
        wait for Clk_period; 
        Features_din <= "0000001001111000";
        wait for Clk_period; 
        Features_din <= "0000001001111000";
        wait for Clk_period; 
        Features_din <= "0000001001111000";
        wait for Clk_period; 
        Features_din <= "0000001001111000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110110111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111111000111000";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "0000000110010001";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "1111111001111100";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000001010100110";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "0000001000000110";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000101000101";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111011101011111";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001000110111";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110011011100";
        wait for Clk_period; 
        Features_din <= "0000001001011011";
        wait for Clk_period; 
        Features_din <= "0000001001011011";
        wait for Clk_period; 
        Features_din <= "0000001001011011";
        wait for Clk_period; 
        Features_din <= "0000001001011011";
        wait for Clk_period; 
        Features_din <= "0000001001011011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110100010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111001000110";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "0000000110001101";
        wait for Clk_period; 
        Features_din <= "0000000011110111";
        wait for Clk_period; 
        Features_din <= "1111111001100001";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000000011110000";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111011110010011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110001111010";
        wait for Clk_period; 
        Features_din <= "0000001001100100";
        wait for Clk_period; 
        Features_din <= "0000001001100100";
        wait for Clk_period; 
        Features_din <= "0000001001100100";
        wait for Clk_period; 
        Features_din <= "0000001001100100";
        wait for Clk_period; 
        Features_din <= "0000001001100100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110111110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111000101001";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "0000000101101011";
        wait for Clk_period; 
        Features_din <= "0000000011111011";
        wait for Clk_period; 
        Features_din <= "1111111001001100";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000011011011";
        wait for Clk_period; 
        Features_din <= "0000000100010011";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000011000010";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111100001001000";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111101101010110";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(3, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111011010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111001010011";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000110000001";
        wait for Clk_period; 
        Features_din <= "0000000011000110";
        wait for Clk_period; 
        Features_din <= "1111111000111000";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000101010010";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111011101011110";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110011011110";
        wait for Clk_period; 
        Features_din <= "0000001001011010";
        wait for Clk_period; 
        Features_din <= "0000001001011010";
        wait for Clk_period; 
        Features_din <= "0000001001011010";
        wait for Clk_period; 
        Features_din <= "0000001001011010";
        wait for Clk_period; 
        Features_din <= "0000001001011010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(6, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110100010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100111111";
        wait for Clk_period; 
        Features_din <= "1111111000100111";
        wait for Clk_period; 
        Features_din <= "1111111110100001";
        wait for Clk_period; 
        Features_din <= "0000000011001111";
        wait for Clk_period; 
        Features_din <= "0000000110010011";
        wait for Clk_period; 
        Features_din <= "0000000100000000";
        wait for Clk_period; 
        Features_din <= "1111111001001110";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000101000001";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "0000000110100011";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "0000000100010111";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000011001000";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111100011000011";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111101010110011";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111001001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111001100000";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "0000000110001110";
        wait for Clk_period; 
        Features_din <= "0000000010101100";
        wait for Clk_period; 
        Features_din <= "1111111000111001";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000011010010";
        wait for Clk_period; 
        Features_din <= "0000000101001101";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000011100101";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "1111011111000110";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110000100000";
        wait for Clk_period; 
        Features_din <= "0000001001101100";
        wait for Clk_period; 
        Features_din <= "0000001001101100";
        wait for Clk_period; 
        Features_din <= "0000001001101100";
        wait for Clk_period; 
        Features_din <= "0000001001101100";
        wait for Clk_period; 
        Features_din <= "0000001001101100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111110101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100100010";
        wait for Clk_period; 
        Features_din <= "1111111001011000";
        wait for Clk_period; 
        Features_din <= "1111111111001010";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000101110111";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "1111111001001110";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000011110111";
        wait for Clk_period; 
        Features_din <= "0000000111000110";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000001000111110";
        wait for Clk_period; 
        Features_din <= "0000000100011001";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000110001110";
        wait for Clk_period; 
        Features_din <= "0000001100010111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "1111111010001011";
        wait for Clk_period; 
        Features_din <= "1111101000111010";
        wait for Clk_period; 
        Features_din <= "0000010010110110";
        wait for Clk_period; 
        Features_din <= "1111110101100110";
        wait for Clk_period; 
        Features_din <= "0000011000110000";
        wait for Clk_period; 
        Features_din <= "1111110101100010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111100011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111000101000";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000101111100";
        wait for Clk_period; 
        Features_din <= "0000000011100001";
        wait for Clk_period; 
        Features_din <= "1111111010000100";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "0000000011111000";
        wait for Clk_period; 
        Features_din <= "0000000100001110";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "1111011101110110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110010101111";
        wait for Clk_period; 
        Features_din <= "0000001001011111";
        wait for Clk_period; 
        Features_din <= "0000001001011111";
        wait for Clk_period; 
        Features_din <= "0000001001011111";
        wait for Clk_period; 
        Features_din <= "0000001001011111";
        wait for Clk_period; 
        Features_din <= "0000001001011111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111110010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111001111000";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000110010110";
        wait for Clk_period; 
        Features_din <= "0000000011000010";
        wait for Clk_period; 
        Features_din <= "1111111001010101";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111011101110001";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110010111001";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111101100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000000110010001";
        wait for Clk_period; 
        Features_din <= "0000000011000101";
        wait for Clk_period; 
        Features_din <= "1111111001000010";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000011101010";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000100000000";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111111010010001";
        wait for Clk_period; 
        Features_din <= "0000000100111001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000001100000010";
        wait for Clk_period; 
        Features_din <= "0000010001111101";
        wait for Clk_period; 
        Features_din <= "1111101111010010";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "1111100100001111";
        wait for Clk_period; 
        Features_din <= "0000000101111000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111001010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100100101";
        wait for Clk_period; 
        Features_din <= "1111111001011000";
        wait for Clk_period; 
        Features_din <= "1111111111000100";
        wait for Clk_period; 
        Features_din <= "0000000011001011";
        wait for Clk_period; 
        Features_din <= "0000000101100000";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "1111111001011111";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "0000000011100001";
        wait for Clk_period; 
        Features_din <= "0000000100110000";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000011000101";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111011110110110";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110000111010";
        wait for Clk_period; 
        Features_din <= "0000001001101001";
        wait for Clk_period; 
        Features_din <= "0000001001101001";
        wait for Clk_period; 
        Features_din <= "0000001001101001";
        wait for Clk_period; 
        Features_din <= "0000001001101001";
        wait for Clk_period; 
        Features_din <= "0000001001101001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111100000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "1111111001010001";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000000110011000";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "1111111000111001";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000101001001";
        wait for Clk_period; 
        Features_din <= "0000000011010000";
        wait for Clk_period; 
        Features_din <= "0000000011110100";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000101110000";
        wait for Clk_period; 
        Features_din <= "0000000100101011";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000011101110";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111100101110110";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111100111100101";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110111111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111001000011";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000000110001100";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "1111111000101110";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000000011101101";
        wait for Clk_period; 
        Features_din <= "0000000011010011";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111011101001010";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111110100000111";
        wait for Clk_period; 
        Features_din <= "0000001001010110";
        wait for Clk_period; 
        Features_din <= "0000001001010110";
        wait for Clk_period; 
        Features_din <= "0000001001010110";
        wait for Clk_period; 
        Features_din <= "0000001001010110";
        wait for Clk_period; 
        Features_din <= "0000001001010110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110101111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111001101111";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000110101111";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "1111111000100001";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000001010101101";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000000100100101";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111100100100100";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001011110000";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111101000111110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111010101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111001011111";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "0000000110100000";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "1111111001000111";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000000011011111";
        wait for Clk_period; 
        Features_din <= "0000000111111010";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "0000000100011101";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111100011010001";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111101010100001";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111010101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111000111001";
        wait for Clk_period; 
        Features_din <= "1111111110110010";
        wait for Clk_period; 
        Features_din <= "0000000100000000";
        wait for Clk_period; 
        Features_din <= "0000000110000010";
        wait for Clk_period; 
        Features_din <= "0000000011111100";
        wait for Clk_period; 
        Features_din <= "1111111001100101";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000011101001";
        wait for Clk_period; 
        Features_din <= "0000001011011100";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111100000010101";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001011001001";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111101110100001";
        wait for Clk_period; 
        Features_din <= "0000001001110101";
        wait for Clk_period; 
        Features_din <= "0000001001110101";
        wait for Clk_period; 
        Features_din <= "0000001001110101";
        wait for Clk_period; 
        Features_din <= "0000001001110101";
        wait for Clk_period; 
        Features_din <= "0000001001110101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(5, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000000001010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100111010";
        wait for Clk_period; 
        Features_din <= "1111111001110010";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000110110010";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111110111111100";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000001100001100";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111100100101110";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001010010100";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111101000110011";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111101001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111001011110";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "0000000110011011";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "1111111001100110";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000011010000";
        wait for Clk_period; 
        Features_din <= "0000000111010001";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000011010101";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000100000001";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "1111101000101101";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "1111100100110100";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111100001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111001011100";
        wait for Clk_period; 
        Features_din <= "1111111110110001";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "0000000101101010";
        wait for Clk_period; 
        Features_din <= "0000000011101100";
        wait for Clk_period; 
        Features_din <= "1111111001011011";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000001000000010";
        wait for Clk_period; 
        Features_din <= "0000000011011101";
        wait for Clk_period; 
        Features_din <= "0000001001001111";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000001000110100";
        wait for Clk_period; 
        Features_din <= "0000000101010100";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111100101101100";
        wait for Clk_period; 
        Features_din <= "0000001100010000";
        wait for Clk_period; 
        Features_din <= "0000001010010011";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111100111110000";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111001001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101000001";
        wait for Clk_period; 
        Features_din <= "1111111001001001";
        wait for Clk_period; 
        Features_din <= "1111111111010110";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000000101110001";
        wait for Clk_period; 
        Features_din <= "0000000011100100";
        wait for Clk_period; 
        Features_din <= "1111111000111010";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000011011010";
        wait for Clk_period; 
        Features_din <= "0000000101100111";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "0000000111101100";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000011001010";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111100001111110";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101100001100";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111010100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111001111010";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "0000000111010101";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "1111111001001100";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000001001010100";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000101000111";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000001010001101";
        wait for Clk_period; 
        Features_din <= "0000001001100110";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000011011100";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000001011111110";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000111100001";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "0000010011110011";
        wait for Clk_period; 
        Features_din <= "0000001011000101";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "1111011101010101";
        wait for Clk_period; 
        Features_din <= "0000000111000111";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111001100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111000110101";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000000101101101";
        wait for Clk_period; 
        Features_din <= "0000000100000011";
        wait for Clk_period; 
        Features_din <= "1111111001101110";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000011110001";
        wait for Clk_period; 
        Features_din <= "0000000011011101";
        wait for Clk_period; 
        Features_din <= "0000001001101011";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "0000000101100100";
        wait for Clk_period; 
        Features_din <= "0000000110111111";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111101011001100";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001100001011";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111100010101110";
        wait for Clk_period; 
        Features_din <= "0000001010000001";
        wait for Clk_period; 
        Features_din <= "0000001010000001";
        wait for Clk_period; 
        Features_din <= "0000001010000001";
        wait for Clk_period; 
        Features_din <= "0000001010000001";
        wait for Clk_period; 
        Features_din <= "0000001010000001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111001111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111111001001001";
        wait for Clk_period; 
        Features_din <= "1111111110101010";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "0000000110001101";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "1111111000110010";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000001000000000";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000001010000000";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000100101110";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111100011011100";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001001100110";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111101010010011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110101010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111001001110";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000000101110011";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "1111111001010001";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000000011101110";
        wait for Clk_period; 
        Features_din <= "0000000101101000";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111011110000101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110010010100";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111101010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101001100";
        wait for Clk_period; 
        Features_din <= "1111111001001111";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "0000000110101101";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "1111111000110100";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111011111101001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101111100110";
        wait for Clk_period; 
        Features_din <= "0000001001110000";
        wait for Clk_period; 
        Features_din <= "0000001001110000";
        wait for Clk_period; 
        Features_din <= "0000001001110000";
        wait for Clk_period; 
        Features_din <= "0000001001110000";
        wait for Clk_period; 
        Features_din <= "0000001001110000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111010011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111110001000";
        wait for Clk_period; 
        Features_din <= "1111111001110011";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "0000000111010110";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "1111111000110101";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111100010000110";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111101100000001";
        wait for Clk_period; 
        Features_din <= "0000001001111111";
        wait for Clk_period; 
        Features_din <= "0000001001111111";
        wait for Clk_period; 
        Features_din <= "0000001001111111";
        wait for Clk_period; 
        Features_din <= "0000001001111111";
        wait for Clk_period; 
        Features_din <= "0000001001111111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111001110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101101000";
        wait for Clk_period; 
        Features_din <= "1111111001110000";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000111001111";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111111000111100";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000111101100";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "0000001001001010";
        wait for Clk_period; 
        Features_din <= "0000000011111011";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "1111101001001111";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000000101000001";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111100100010110";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111111000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111001011000";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "0000000011000001";
        wait for Clk_period; 
        Features_din <= "0000000101011010";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "1111111001101110";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000000011100111";
        wait for Clk_period; 
        Features_din <= "0000000111100011";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111100000011100";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101110010110";
        wait for Clk_period; 
        Features_din <= "0000001001110110";
        wait for Clk_period; 
        Features_din <= "0000001001110110";
        wait for Clk_period; 
        Features_din <= "0000001001110110";
        wait for Clk_period; 
        Features_din <= "0000001001110110";
        wait for Clk_period; 
        Features_din <= "0000001001110110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111011100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101011101";
        wait for Clk_period; 
        Features_din <= "1111111001000001";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "0000000011001001";
        wait for Clk_period; 
        Features_din <= "0000000110010011";
        wait for Clk_period; 
        Features_din <= "0000000011000000";
        wait for Clk_period; 
        Features_din <= "1111111001011011";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000011101110";
        wait for Clk_period; 
        Features_din <= "0000000100001011";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111011110100010";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110001011110";
        wait for Clk_period; 
        Features_din <= "0000001001100110";
        wait for Clk_period; 
        Features_din <= "0000001001100110";
        wait for Clk_period; 
        Features_din <= "0000001001100110";
        wait for Clk_period; 
        Features_din <= "0000001001100110";
        wait for Clk_period; 
        Features_din <= "0000001001100110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110100101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111001000110";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000000101111001";
        wait for Clk_period; 
        Features_din <= "0000000011000100";
        wait for Clk_period; 
        Features_din <= "1111111001011000";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000111111111";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "0000001100101101";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000010111110";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111011111100110";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000000101100010";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101111101011";
        wait for Clk_period; 
        Features_din <= "0000001001110000";
        wait for Clk_period; 
        Features_din <= "0000001001110000";
        wait for Clk_period; 
        Features_din <= "0000001001110000";
        wait for Clk_period; 
        Features_din <= "0000001001110000";
        wait for Clk_period; 
        Features_din <= "0000001001110000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111010110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101000010";
        wait for Clk_period; 
        Features_din <= "1111111001111101";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000110011000";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "1111111000111100";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000001001000111";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "0000001011110111";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000001001101101";
        wait for Clk_period; 
        Features_din <= "0000000100110011";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000010110010";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "1111101000001100";
        wait for Clk_period; 
        Features_din <= "0000001011110010";
        wait for Clk_period; 
        Features_din <= "0000000101101011";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111100101010010";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111011000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111001010010";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "0000000010110010";
        wait for Clk_period; 
        Features_din <= "0000000101010101";
        wait for Clk_period; 
        Features_din <= "0000000010111111";
        wait for Clk_period; 
        Features_din <= "1111111001100111";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000011100110";
        wait for Clk_period; 
        Features_din <= "0000001000001101";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000000011011010";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000010111000";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111011111100001";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111101111110010";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111011010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111000111101";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "0000000110011100";
        wait for Clk_period; 
        Features_din <= "0000000011010111";
        wait for Clk_period; 
        Features_din <= "1111111000011111";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000001001001100";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000110011011";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "0000000111100100";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000011110110";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111100010111011";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001011011011";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111101010111100";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111001000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111000100111";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "0000000011000110";
        wait for Clk_period; 
        Features_din <= "0000000110001011";
        wait for Clk_period; 
        Features_din <= "0000000011010000";
        wait for Clk_period; 
        Features_din <= "1111111001101010";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000100000000";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111011010111101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111001100011";
        wait for Clk_period; 
        Features_din <= "0000001000101101";
        wait for Clk_period; 
        Features_din <= "0000001000101101";
        wait for Clk_period; 
        Features_din <= "0000001000101101";
        wait for Clk_period; 
        Features_din <= "0000001000101101";
        wait for Clk_period; 
        Features_din <= "0000001000101101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110110001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111000000101";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "0000000100000101";
        wait for Clk_period; 
        Features_din <= "0000000100111000";
        wait for Clk_period; 
        Features_din <= "0000000100101101";
        wait for Clk_period; 
        Features_din <= "1111111001111100";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "0000000011111001";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111011110110011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110001000001";
        wait for Clk_period; 
        Features_din <= "0000001001101001";
        wait for Clk_period; 
        Features_din <= "0000001001101001";
        wait for Clk_period; 
        Features_din <= "0000001001101001";
        wait for Clk_period; 
        Features_din <= "0000001001101001";
        wait for Clk_period; 
        Features_din <= "0000001001101001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111011100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100101101";
        wait for Clk_period; 
        Features_din <= "1111111001000101";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000000101101010";
        wait for Clk_period; 
        Features_din <= "0000000011011001";
        wait for Clk_period; 
        Features_din <= "1111111001000011";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000001001100000";
        wait for Clk_period; 
        Features_din <= "0000000011101010";
        wait for Clk_period; 
        Features_din <= "0000001000111000";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000110010100";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111011111011111";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001001010101";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111101111110111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111011011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "1111111000111000";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "0000000110101011";
        wait for Clk_period; 
        Features_din <= "0000000011011101";
        wait for Clk_period; 
        Features_din <= "1111111001010110";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000011110010";
        wait for Clk_period; 
        Features_din <= "0000000111010111";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111100010100100";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101011011001";
        wait for Clk_period; 
        Features_din <= "0000001010000001";
        wait for Clk_period; 
        Features_din <= "0000001010000001";
        wait for Clk_period; 
        Features_din <= "0000001010000001";
        wait for Clk_period; 
        Features_din <= "0000001010000001";
        wait for Clk_period; 
        Features_din <= "0000001010000001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111010010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101011011";
        wait for Clk_period; 
        Features_din <= "1111111001110001";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000000111111010";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111111001010010";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000001011010001";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "0000001011010100";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000001000111101";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111100101101011";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111100111110001";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111001010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111001100100";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000110001010";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "1111111001101001";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "0000000101011101";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111011101011000";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110011101011";
        wait for Clk_period; 
        Features_din <= "0000001001011001";
        wait for Clk_period; 
        Features_din <= "0000001001011001";
        wait for Clk_period; 
        Features_din <= "0000001001011001";
        wait for Clk_period; 
        Features_din <= "0000001001011001";
        wait for Clk_period; 
        Features_din <= "0000001001011001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110111111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111000110111";
        wait for Clk_period; 
        Features_din <= "1111111111011111";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "0000000110010110";
        wait for Clk_period; 
        Features_din <= "0000000011011001";
        wait for Clk_period; 
        Features_din <= "1111111001001010";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000101000001";
        wait for Clk_period; 
        Features_din <= "0000000011100011";
        wait for Clk_period; 
        Features_din <= "0000000110101011";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000000011111000";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000010110011";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111011111010100";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111110000001001";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(3, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110111110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111110001001";
        wait for Clk_period; 
        Features_din <= "1111111001010001";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000111010101";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "1111111001000100";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000001010001100";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000001100010101";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111011111010100";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000000010111000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110000001001";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111000011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100111101";
        wait for Clk_period; 
        Features_din <= "1111111001100100";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000110001111";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "1111111001010101";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000000110101101";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000001001011000";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000010101101";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "1111100000101100";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000000011010101";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101101111111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111000001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111000101001";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "0000000110010010";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "0000000011011100";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000011000000";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111011110101000";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110001010100";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111011101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111111000101001";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "0000000101110101";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "1111111001101011";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000011111010";
        wait for Clk_period; 
        Features_din <= "0000000011011011";
        wait for Clk_period; 
        Features_din <= "0000000100101010";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "1111011110000100";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110010010100";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111110101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100101100";
        wait for Clk_period; 
        Features_din <= "1111111001010001";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "0000000110010111";
        wait for Clk_period; 
        Features_din <= "0000000011001001";
        wait for Clk_period; 
        Features_din <= "1111111001101000";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000101011100";
        wait for Clk_period; 
        Features_din <= "0000000011000001";
        wait for Clk_period; 
        Features_din <= "0000000101111011";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000010101100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111011101010010";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110011110110";
        wait for Clk_period; 
        Features_din <= "0000001001011000";
        wait for Clk_period; 
        Features_din <= "0000001001011000";
        wait for Clk_period; 
        Features_din <= "0000001001011000";
        wait for Clk_period; 
        Features_din <= "0000001001011000";
        wait for Clk_period; 
        Features_din <= "0000001001011000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111010100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "1111111000011000";
        wait for Clk_period; 
        Features_din <= "1111111110001110";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000000110000011";
        wait for Clk_period; 
        Features_din <= "0000000011110000";
        wait for Clk_period; 
        Features_din <= "1111111010001011";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000000011100010";
        wait for Clk_period; 
        Features_din <= "0000000101101101";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000000101000000";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "1111100000100100";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101110001010";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111110011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111111000111101";
        wait for Clk_period; 
        Features_din <= "1111111111010100";
        wait for Clk_period; 
        Features_din <= "0000000010101100";
        wait for Clk_period; 
        Features_din <= "0000000110001111";
        wait for Clk_period; 
        Features_din <= "0000000011010011";
        wait for Clk_period; 
        Features_din <= "1111111001000110";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000011011100";
        wait for Clk_period; 
        Features_din <= "0000001000010101";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000001001000001";
        wait for Clk_period; 
        Features_din <= "0000000101001000";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000011010010";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111100111110010";
        wait for Clk_period; 
        Features_din <= "0000001100001100";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111100101101010";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(5, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111000001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111000101111";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "0000000010110011";
        wait for Clk_period; 
        Features_din <= "0000000101101100";
        wait for Clk_period; 
        Features_din <= "0000000011010101";
        wait for Clk_period; 
        Features_din <= "1111111001010000";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "0000000011101011";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111011100110101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110100110100";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110101000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111001001000";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "0000000110011011";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "1111111001010110";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "0000000110000010";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "0000000100000011";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000011001110";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111011100110001";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110100111100";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111000001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111001001101";
        wait for Clk_period; 
        Features_din <= "1111111111001000";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000110001111";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "1111111001101110";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000100001001";
        wait for Clk_period; 
        Features_din <= "0000000011011100";
        wait for Clk_period; 
        Features_din <= "0000000100000100";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000011000101";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111011111000011";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110000100101";
        wait for Clk_period; 
        Features_din <= "0000001001101011";
        wait for Clk_period; 
        Features_din <= "0000001001101011";
        wait for Clk_period; 
        Features_din <= "0000001001101011";
        wait for Clk_period; 
        Features_din <= "0000001001101011";
        wait for Clk_period; 
        Features_din <= "0000001001101011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111000101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100101001";
        wait for Clk_period; 
        Features_din <= "1111111001101111";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "0000000110001110";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "1111111000101010";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111011100100101";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110101010111";
        wait for Clk_period; 
        Features_din <= "0000001001001110";
        wait for Clk_period; 
        Features_din <= "0000001001001110";
        wait for Clk_period; 
        Features_din <= "0000001001001110";
        wait for Clk_period; 
        Features_din <= "0000001001001110";
        wait for Clk_period; 
        Features_din <= "0000001001001110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111101010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111001001110";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "0000000110010001";
        wait for Clk_period; 
        Features_din <= "0000000011001101";
        wait for Clk_period; 
        Features_din <= "1111111001010100";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000011100001";
        wait for Clk_period; 
        Features_din <= "0000000101110100";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000101000101";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010111100";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111100011010010";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111101010100000";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110101000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111000110110";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "0000000010111111";
        wait for Clk_period; 
        Features_din <= "0000000100111010";
        wait for Clk_period; 
        Features_din <= "0000000100000100";
        wait for Clk_period; 
        Features_din <= "1111111001110001";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "0000000011101111";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111011101100110";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110011001111";
        wait for Clk_period; 
        Features_din <= "0000001001011100";
        wait for Clk_period; 
        Features_din <= "0000001001011100";
        wait for Clk_period; 
        Features_din <= "0000001001011100";
        wait for Clk_period; 
        Features_din <= "0000001001011100";
        wait for Clk_period; 
        Features_din <= "0000001001011100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111000000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111001010011";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "0000000101111011";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "1111111001101000";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000011100111";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111011100010111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111110101110111";
        wait for Clk_period; 
        Features_din <= "0000001001001010";
        wait for Clk_period; 
        Features_din <= "0000001001001010";
        wait for Clk_period; 
        Features_din <= "0000001001001010";
        wait for Clk_period; 
        Features_din <= "0000001001001010";
        wait for Clk_period; 
        Features_din <= "0000001001001010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111000011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100100100";
        wait for Clk_period; 
        Features_din <= "1111111000010011";
        wait for Clk_period; 
        Features_din <= "1111111110110111";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "0000000101101011";
        wait for Clk_period; 
        Features_din <= "0000000011011010";
        wait for Clk_period; 
        Features_din <= "1111111001101100";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "0000000011011110";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000011000010";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111011011111010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110110111101";
        wait for Clk_period; 
        Features_din <= "0000001001000010";
        wait for Clk_period; 
        Features_din <= "0000001001000010";
        wait for Clk_period; 
        Features_din <= "0000001001000010";
        wait for Clk_period; 
        Features_din <= "0000001001000010";
        wait for Clk_period; 
        Features_din <= "0000001001000010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(5, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111101001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111001100011";
        wait for Clk_period; 
        Features_din <= "1111111110111101";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000110001101";
        wait for Clk_period; 
        Features_din <= "0000000011010010";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000100010000";
        wait for Clk_period; 
        Features_din <= "0000000011100100";
        wait for Clk_period; 
        Features_din <= "0000001001001111";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000100100110";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111100001011000";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001100010111";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111101101000000";
        wait for Clk_period; 
        Features_din <= "0000001001111011";
        wait for Clk_period; 
        Features_din <= "0000001001111011";
        wait for Clk_period; 
        Features_din <= "0000001001111011";
        wait for Clk_period; 
        Features_din <= "0000001001111011";
        wait for Clk_period; 
        Features_din <= "0000001001111011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111011110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111001111111";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "0000000111011010";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "1111111000101010";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000110111100";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "1111101000110011";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "1111100100101110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001000110001";
        wait for Clk_period; 
        Features_din <= "0000001100010111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000101000111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110101001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "1111111001001010";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "0000000110111001";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "1111111001000001";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000010111111";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111011101100100";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110011010011";
        wait for Clk_period; 
        Features_din <= "0000001001011011";
        wait for Clk_period; 
        Features_din <= "0000001001011011";
        wait for Clk_period; 
        Features_din <= "0000001001011011";
        wait for Clk_period; 
        Features_din <= "0000001001011011";
        wait for Clk_period; 
        Features_din <= "0000001001011011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111010010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111111001001010";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000000110010100";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "1111111000111001";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "1111011110000011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110010011000";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111100111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100110101";
        wait for Clk_period; 
        Features_din <= "1111111001100001";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000000110001111";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "1111111001001100";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000110000101";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000110000100";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000000010111110";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111100101100001";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000000110111000";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111100111111011";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(3, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111010001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100110111";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000000110110101";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "1111111000011010";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111100001001101";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101101001111";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111001101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111001011010";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000000110000101";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "1111111001100101";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000011100111";
        wait for Clk_period; 
        Features_din <= "0000000100010001";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111011111110011";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101111010101";
        wait for Clk_period; 
        Features_din <= "0000001001110001";
        wait for Clk_period; 
        Features_din <= "0000001001110001";
        wait for Clk_period; 
        Features_din <= "0000001001110001";
        wait for Clk_period; 
        Features_din <= "0000001001110001";
        wait for Clk_period; 
        Features_din <= "0000001001110001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111010111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100110100";
        wait for Clk_period; 
        Features_din <= "1111111000110110";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "0000000011001111";
        wait for Clk_period; 
        Features_din <= "0000000101010101";
        wait for Clk_period; 
        Features_din <= "0000000100010111";
        wait for Clk_period; 
        Features_din <= "1111111001010110";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000011111000";
        wait for Clk_period; 
        Features_din <= "0000000011011100";
        wait for Clk_period; 
        Features_din <= "0000001011111110";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "0000000110000110";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111100111111010";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001001111001";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111100101100010";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111011011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111010011011";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000110011100";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "1111111000100000";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "0000000110000001";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "0000000011100000";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000011001100";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "1111100011101010";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111101010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111110000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111111001011110";
        wait for Clk_period; 
        Features_din <= "1111111111100000";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000000110010100";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000001000101011";
        wait for Clk_period; 
        Features_din <= "0000000011100010";
        wait for Clk_period; 
        Features_din <= "0000000111110111";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "0000000101001010";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111100000011100";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001010111010";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111101110010111";
        wait for Clk_period; 
        Features_din <= "0000001001110110";
        wait for Clk_period; 
        Features_din <= "0000001001110110";
        wait for Clk_period; 
        Features_din <= "0000001001110110";
        wait for Clk_period; 
        Features_din <= "0000001001110110";
        wait for Clk_period; 
        Features_din <= "0000001001110110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111010011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "1111111001010101";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "0000000010101101";
        wait for Clk_period; 
        Features_din <= "0000000110011001";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "1111111000100010";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111011110001100";
        wait for Clk_period; 
        Features_din <= "0000001000111100";
        wait for Clk_period; 
        Features_din <= "0000000010111100";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110010000111";
        wait for Clk_period; 
        Features_din <= "0000001001100011";
        wait for Clk_period; 
        Features_din <= "0000001001100011";
        wait for Clk_period; 
        Features_din <= "0000001001100011";
        wait for Clk_period; 
        Features_din <= "0000001001100011";
        wait for Clk_period; 
        Features_din <= "0000001001100011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111100001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111111001100011";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "0000000110001010";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "1111111001000101";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000010111110";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111011110000110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110010010001";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111010011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100011010";
        wait for Clk_period; 
        Features_din <= "1111111000100101";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "0000000110000001";
        wait for Clk_period; 
        Features_din <= "0000000011010001";
        wait for Clk_period; 
        Features_din <= "1111111001100111";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000110000101";
        wait for Clk_period; 
        Features_din <= "0000000011100011";
        wait for Clk_period; 
        Features_din <= "0000001001111101";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000001000100000";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000010101101";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111100010011000";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001010111101";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111101011101000";
        wait for Clk_period; 
        Features_din <= "0000001010000000";
        wait for Clk_period; 
        Features_din <= "0000001010000000";
        wait for Clk_period; 
        Features_din <= "0000001010000000";
        wait for Clk_period; 
        Features_din <= "0000001010000000";
        wait for Clk_period; 
        Features_din <= "0000001010000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111011111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101100110";
        wait for Clk_period; 
        Features_din <= "1111111001100000";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000000110110110";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "1111111000110001";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000001011010111";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000001010111010";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000000111110001";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111100011011101";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111101010010010";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111000001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101010100";
        wait for Clk_period; 
        Features_din <= "1111111001010110";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "0000000011001000";
        wait for Clk_period; 
        Features_din <= "0000000101100111";
        wait for Clk_period; 
        Features_din <= "0000000011101011";
        wait for Clk_period; 
        Features_din <= "1111111001010010";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000011101010";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111011101110101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110010110001";
        wait for Clk_period; 
        Features_din <= "0000001001011111";
        wait for Clk_period; 
        Features_din <= "0000001001011111";
        wait for Clk_period; 
        Features_din <= "0000001001011111";
        wait for Clk_period; 
        Features_din <= "0000001001011111";
        wait for Clk_period; 
        Features_din <= "0000001001011111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111010110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111000111001";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "0000000110010100";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "1111111001100101";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000001010011100";
        wait for Clk_period; 
        Features_din <= "0000000011101011";
        wait for Clk_period; 
        Features_din <= "0000000111001011";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000000110011010";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111011110100011";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001001110010";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110001011100";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111100101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111111001111000";
        wait for Clk_period; 
        Features_din <= "1111111111010101";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "0000000110101001";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "1111111001000111";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000000011110001";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000001000111101";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111100010010110";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000000110000110";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101011101011";
        wait for Clk_period; 
        Features_din <= "0000001010000000";
        wait for Clk_period; 
        Features_din <= "0000001010000000";
        wait for Clk_period; 
        Features_din <= "0000001010000000";
        wait for Clk_period; 
        Features_din <= "0000001010000000";
        wait for Clk_period; 
        Features_din <= "0000001010000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111001111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101000011";
        wait for Clk_period; 
        Features_din <= "1111111000111001";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "0000000010110010";
        wait for Clk_period; 
        Features_din <= "0000000101111111";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "1111111001011010";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000011000000";
        wait for Clk_period; 
        Features_din <= "0000000011100001";
        wait for Clk_period; 
        Features_din <= "0000000111100011";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000011000010";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111011111010100";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111110000001001";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111110010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100111100";
        wait for Clk_period; 
        Features_din <= "1111111000110010";
        wait for Clk_period; 
        Features_din <= "1111111111010111";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000000110010101";
        wait for Clk_period; 
        Features_din <= "0000000010111000";
        wait for Clk_period; 
        Features_din <= "1111111001011100";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000111111100";
        wait for Clk_period; 
        Features_din <= "0000000011110001";
        wait for Clk_period; 
        Features_din <= "0000000111011010";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000100010100";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111100000000000";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001011110000";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111101111000010";
        wait for Clk_period; 
        Features_din <= "0000001001110011";
        wait for Clk_period; 
        Features_din <= "0000001001110011";
        wait for Clk_period; 
        Features_din <= "0000001001110011";
        wait for Clk_period; 
        Features_din <= "0000001001110011";
        wait for Clk_period; 
        Features_din <= "0000001001110011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110111000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111111000110101";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000000110010110";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "1111111000010011";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000001100001101";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000100010100";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111100011101000";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001010000001";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111101010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111011011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100001110";
        wait for Clk_period; 
        Features_din <= "1111111001010101";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "0000000101110101";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "1111111001110100";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000011000101";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111011101110010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110010111000";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(5, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111011011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100100001";
        wait for Clk_period; 
        Features_din <= "1111111001000101";
        wait for Clk_period; 
        Features_din <= "1111111111000101";
        wait for Clk_period; 
        Features_din <= "0000000011001001";
        wait for Clk_period; 
        Features_din <= "0000000101111011";
        wait for Clk_period; 
        Features_din <= "0000000011110011";
        wait for Clk_period; 
        Features_din <= "1111111001101000";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000011100001";
        wait for Clk_period; 
        Features_din <= "0000000010111111";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111100001100001";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111101100110011";
        wait for Clk_period; 
        Features_din <= "0000001001111100";
        wait for Clk_period; 
        Features_din <= "0000001001111100";
        wait for Clk_period; 
        Features_din <= "0000001001111100";
        wait for Clk_period; 
        Features_din <= "0000001001111100";
        wait for Clk_period; 
        Features_din <= "0000001001111100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111011011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100011001";
        wait for Clk_period; 
        Features_din <= "1111111000101010";
        wait for Clk_period; 
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000000110010000";
        wait for Clk_period; 
        Features_din <= "0000000011100100";
        wait for Clk_period; 
        Features_din <= "1111111001011101";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "0000001000000001";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000110101000";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111011110011010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000000011011010";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110001101100";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111001011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100110110";
        wait for Clk_period; 
        Features_din <= "1111111000111111";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "0000000110000011";
        wait for Clk_period; 
        Features_din <= "0000000011000101";
        wait for Clk_period; 
        Features_din <= "1111111001001101";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000111100100";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "0000001001001111";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000011010001";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111011111010111";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001010101010";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111110000000011";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111110011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "1111111001110111";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "0000000110101110";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "1111111001000100";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000111100000";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000001000111010";
        wait for Clk_period; 
        Features_din <= "0000000110011110";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111101010001101";
        wait for Clk_period; 
        Features_din <= "0000001011100111";
        wait for Clk_period; 
        Features_din <= "0000000101010011";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111100011100001";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(6, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110011110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111111000011110";
        wait for Clk_period; 
        Features_din <= "1111111111110001";
        wait for Clk_period; 
        Features_din <= "0000000011001010";
        wait for Clk_period; 
        Features_din <= "0000000111100011";
        wait for Clk_period; 
        Features_din <= "0000000011011001";
        wait for Clk_period; 
        Features_din <= "1111111000011000";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000001100110010";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000100111011";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000001010101000";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000011110000";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111100011001010";
        wait for Clk_period; 
        Features_din <= "0000001011111101";
        wait for Clk_period; 
        Features_din <= "0000001000010010";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111101010101001";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110110000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100100111";
        wait for Clk_period; 
        Features_din <= "1111111000010001";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "0000000101010111";
        wait for Clk_period; 
        Features_din <= "0000000100001100";
        wait for Clk_period; 
        Features_din <= "1111111001011110";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "0000000011101001";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000010110010";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "1111011110100110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110001010111";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111010000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "1111111001100101";
        wait for Clk_period; 
        Features_din <= "1111111111100111";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000110001001";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "1111111000111011";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000010101101";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111100001111001";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111101100010010";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111011101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "1111111001010100";
        wait for Clk_period; 
        Features_din <= "1111111111001101";
        wait for Clk_period; 
        Features_din <= "0000000011000111";
        wait for Clk_period; 
        Features_din <= "0000000101111100";
        wait for Clk_period; 
        Features_din <= "0000000010101100";
        wait for Clk_period; 
        Features_din <= "1111111001011111";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000111111101";
        wait for Clk_period; 
        Features_din <= "0000000011011001";
        wait for Clk_period; 
        Features_din <= "0000001001010101";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000001000001100";
        wait for Clk_period; 
        Features_din <= "0000000011111000";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010110010";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111100100001010";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001010010010";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111101001011101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111011100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101101010";
        wait for Clk_period; 
        Features_din <= "1111111010000110";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000000111011010";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "1111111000000001";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "1111011111011111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101111110101";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111101100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100011101";
        wait for Clk_period; 
        Features_din <= "1111111001100011";
        wait for Clk_period; 
        Features_din <= "1111111111011001";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000101000000";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "1111111001000110";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000011101111";
        wait for Clk_period; 
        Features_din <= "0000000110110000";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000100011100";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000100001101";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111101001010110";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "1111100100010000";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111110111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101000100";
        wait for Clk_period; 
        Features_din <= "1111111001101001";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000111010011";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111111001011101";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000001100011010";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000001000101111";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "0000000101111010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111100001000001";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000000101000110";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101101011111";
        wait for Clk_period; 
        Features_din <= "0000001001111001";
        wait for Clk_period; 
        Features_din <= "0000001001111001";
        wait for Clk_period; 
        Features_din <= "0000001001111001";
        wait for Clk_period; 
        Features_din <= "0000001001111001";
        wait for Clk_period; 
        Features_din <= "0000001001111001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111000101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100010100";
        wait for Clk_period; 
        Features_din <= "1111111001011110";
        wait for Clk_period; 
        Features_din <= "1111111111010011";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "0000000101110000";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "1111111001100110";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000011100000";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000011000111";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111011101000100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110100010101";
        wait for Clk_period; 
        Features_din <= "0000001001010101";
        wait for Clk_period; 
        Features_din <= "0000001001010101";
        wait for Clk_period; 
        Features_din <= "0000001001010101";
        wait for Clk_period; 
        Features_din <= "0000001001010101";
        wait for Clk_period; 
        Features_din <= "0000001001010101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(5, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110111000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101001010";
        wait for Clk_period; 
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000111000100";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "1111111000111110";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000101111001";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000001100010101";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000100100110";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "1111100011111111";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001000010101";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111101001101010";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111000111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "1111111001000100";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "0000000011000000";
        wait for Clk_period; 
        Features_din <= "0000000110000110";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "1111111001000001";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000000011100000";
        wait for Clk_period; 
        Features_din <= "0000001010001010";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000000100010100";
        wait for Clk_period; 
        Features_din <= "0000000011011000";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111100001101001";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001100000111";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111101100101000";
        wait for Clk_period; 
        Features_din <= "0000001001111101";
        wait for Clk_period; 
        Features_din <= "0000001001111101";
        wait for Clk_period; 
        Features_din <= "0000001001111101";
        wait for Clk_period; 
        Features_din <= "0000001001111101";
        wait for Clk_period; 
        Features_din <= "0000001001111101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(6, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111010001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "1111111001000000";
        wait for Clk_period; 
        Features_din <= "1111111111011110";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "0000000101100101";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "1111111001111011";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000001100001010";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000000101000000";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "0000001010110110";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000100010110";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "1111100000101100";
        wait for Clk_period; 
        Features_din <= "0000001011101100";
        wait for Clk_period; 
        Features_din <= "0000001001001000";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101101111111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111010001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101010010";
        wait for Clk_period; 
        Features_din <= "1111111001010101";
        wait for Clk_period; 
        Features_din <= "1111111111101101";
        wait for Clk_period; 
        Features_din <= "0000000011010000";
        wait for Clk_period; 
        Features_din <= "0000000101111100";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "1111111001100001";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000101101000";
        wait for Clk_period; 
        Features_din <= "0000000011110100";
        wait for Clk_period; 
        Features_din <= "0000001000111001";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000000011011000";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111011111000011";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001100000011";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110000100101";
        wait for Clk_period; 
        Features_din <= "0000001001101011";
        wait for Clk_period; 
        Features_din <= "0000001001101011";
        wait for Clk_period; 
        Features_din <= "0000001001101011";
        wait for Clk_period; 
        Features_din <= "0000001001101011";
        wait for Clk_period; 
        Features_din <= "0000001001101011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110111010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "0000000010101101";
        wait for Clk_period; 
        Features_din <= "0000000101111101";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "1111111001001110";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000011101001";
        wait for Clk_period; 
        Features_din <= "0000000011001000";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "1111011011111001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110111000000";
        wait for Clk_period; 
        Features_din <= "0000001001000001";
        wait for Clk_period; 
        Features_din <= "0000001001000001";
        wait for Clk_period; 
        Features_din <= "0000001001000001";
        wait for Clk_period; 
        Features_din <= "0000001001000001";
        wait for Clk_period; 
        Features_din <= "0000001001000001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111101101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111111001001000";
        wait for Clk_period; 
        Features_din <= "1111111111010010";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "0000000101110110";
        wait for Clk_period; 
        Features_din <= "0000000011011111";
        wait for Clk_period; 
        Features_din <= "1111111001000001";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000011101101";
        wait for Clk_period; 
        Features_din <= "0000000110111100";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000000110101101";
        wait for Clk_period; 
        Features_din <= "0000000100011010";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111100101100010";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111100111111010";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(5, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110110001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111111000011110";
        wait for Clk_period; 
        Features_din <= "1111111111010000";
        wait for Clk_period; 
        Features_din <= "0000000010111101";
        wait for Clk_period; 
        Features_din <= "0000000110010000";
        wait for Clk_period; 
        Features_din <= "0000000011010110";
        wait for Clk_period; 
        Features_din <= "1111111001111000";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000011011011";
        wait for Clk_period; 
        Features_din <= "0000000110101011";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "0000000011010110";
        wait for Clk_period; 
        Features_din <= "0000000011010101";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "1111100101111100";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111100111011111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111111000011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100111110";
        wait for Clk_period; 
        Features_din <= "1111111001110010";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "0000000101100110";
        wait for Clk_period; 
        Features_din <= "0000000011010101";
        wait for Clk_period; 
        Features_din <= "1111111001010110";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "0000000100001101";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000010111111";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111100000101011";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111101110000000";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
            wait;
    end process;
end;
