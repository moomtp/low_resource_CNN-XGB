

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.types.all;

entity image_test is
    generic(TREE_RAM_BITS: positive := 14;
            NUM_CLASSES:   positive := 7;
            NUM_FEATURES:  positive := 35);
end image_test;

architecture behavior of image_test is
    
    component image
        generic(TREE_RAM_BITS: positive;
                NUM_CLASSES:   positive;
                NUM_FEATURES:  positive);
        port(-- Control signals
             Clk:   in std_logic;
             Reset: in std_logic;
             
             -- Inputs for the nodes reception (trees)
             Load_trees: in std_logic;
             Valid_node: in std_logic;
             Addr:       in std_logic_vector(TREE_RAM_BITS - 1  downto 0);
             Trees_din:  in std_logic_vector(31 downto 0);
             
             -- Inputs for the features reception (pixels)
             Load_features: in std_logic;
             Valid_feature: in std_logic;
             Features_din:  in std_logic_vector(15 downto 0);
             Last_feature:  in std_logic;
             
             -- Output signals
             --     Finish:     finish (also 'ready') signal
             --     Dout:       the selected class
             --     Greater:    the value of the selected class prediction
             --     Curr_state: the current state
             Finish:     out std_logic;
             Dout:       out std_logic_vector(log_2(NUM_CLASSES) - 1 downto 0);
             greater:    out std_logic_vector(31 downto 0);
             curr_state: out std_logic_vector(2 downto 0));
    end component;
    
    component counter is
        generic(BITS: natural);
        port(Clk:   in  std_logic;
             Reset: in  std_logic;
             Count: in  std_logic;
             Dout:  out std_logic_vector (BITS - 1 downto 0));
    end component;
    
    -- Inputs
    signal Clk:           std_logic := '0';
    signal Reset:         std_logic := '0';
    signal Load_trees:    std_logic := '0';
    signal Valid_node:    std_logic := '0';
    signal Addr:          std_logic_vector(TREE_RAM_BITS - 1 downto
                                           0) := (others => '0');
    signal Trees_din:     std_logic_vector(31 downto 0) := (others => '0');
    signal Load_features: std_logic := '0';
    signal Valid_feature: std_logic := '0';
    signal Features_din:  std_logic_vector(15 downto 0) := (others => '0');
    signal last_feature:  std_logic := '0';
    
    -- Outputs
    signal Finish:     std_logic;
    signal Dout:       std_logic_vector(log_2(NUM_CLASSES) - 1 downto 0);
    signal greater:    std_logic_vector(31 downto 0);
    signal curr_state: std_logic_vector(2 downto 0);
    
    -- Clock period definition
    constant Clk_period : time := 10 ns;
    
    -- Counter signals
    signal pc_count, hc_count: std_logic := '0';
    signal pixels, hits: std_logic_vector(15 downto 0) := (others => '0');
    
    -- Label signal
    signal class_label: std_logic_vector(log_2(NUM_CLASSES) - 1 downto 0);

begin
    
    -- Instantiate the Unit Under Test (UUT)
    uut: image
        generic map(TREE_RAM_BITS => TREE_RAM_BITS,
                    NUM_CLASSES   => NUM_CLASSES,
                    NUM_FEATURES  => NUM_FEATURES)
        port map(Clk           => Clk,
                 Reset         => Reset,
                 Load_trees    => Load_trees,
                 Valid_node    => Valid_node,
                 Addr          => Addr,
                 Trees_din     => Trees_din,
                 Load_features => Load_features,
                 Valid_feature => Valid_feature,
                 Features_din  => Features_din,
                 Last_feature  => Last_feature,
                 Finish        => Finish,
                 Dout          => Dout,
                 greater       => greater,
                 curr_state    => curr_state);
    
    -- To count the pixels
    pixel_counter: counter
        generic map(BITS => 16)
        port map(Clk   => Clk, 
                 Reset => Reset,
                 Count => pc_count,
                 Dout  => pixels);
    
    -- To count the hits
    hit_counter: counter
        generic map(BITS => 16)
        port map(Clk   => Clk, 
                 Reset => Reset,
                 Count => hc_count,
                 Dout  => hits);
    
    -- Clock process definition
    Clk_process: process
    begin
        Clk <= '0';
        wait for Clk_period/2;
        Clk <= '1';
        wait for Clk_period/2;
    end process;
    
    -- Stimulus process
    stim_proc: process
    begin
        
        Reset <= '1';
        
        -- hold reset state for 100 ns.
        wait for 100 ns;
        
        Reset <= '0';
        
        wait for Clk_period*10;
        


        
        -- LOAD TREES
        -----------------------------------------------------------------------
        
        -- Load and valid trees flags
        Load_trees <= '1';
        Valid_node <= '1';

        -- Class  0
        -----------
		Addr <=  "00000000000000";
		Trees_din <= x"050b0748";
		wait for Clk_period;
		Addr <=  "00000000000001";
		Trees_din <= x"0508551c";
		wait for Clk_period;
		Addr <=  "00000000000010";
		Trees_din <= x"0506f70c";
		wait for Clk_period;
		Addr <=  "00000000000011";
		Trees_din <= x"20000e04";
		wait for Clk_period;
		Addr <=  "00000000000100";
		Trees_din <= x"ff4d00ed";
		wait for Clk_period;
		Addr <=  "00000000000101";
		Trees_din <= x"03fe1f04";
		wait for Clk_period;
		Addr <=  "00000000000110";
		Trees_din <= x"002700ed";
		wait for Clk_period;
		Addr <=  "00000000000111";
		Trees_din <= x"ff7100ed";
		wait for Clk_period;
		Addr <=  "00000000001000";
		Trees_din <= x"04fd7604";
		wait for Clk_period;
		Addr <=  "00000000001001";
		Trees_din <= x"010400ed";
		wait for Clk_period;
		Addr <=  "00000000001010";
		Trees_din <= x"1c005108";
		wait for Clk_period;
		Addr <=  "00000000001011";
		Trees_din <= x"0bf98004";
		wait for Clk_period;
		Addr <=  "00000000001100";
		Trees_din <= x"ffd000ed";
		wait for Clk_period;
		Addr <=  "00000000001101";
		Trees_din <= x"ff5100ed";
		wait for Clk_period;
		Addr <=  "00000000001110";
		Trees_din <= x"008e00ed";
		wait for Clk_period;
		Addr <=  "00000000001111";
		Trees_din <= x"03fc8810";
		wait for Clk_period;
		Addr <=  "00000000010000";
		Trees_din <= x"0a008c08";
		wait for Clk_period;
		Addr <=  "00000000010001";
		Trees_din <= x"03fb1e04";
		wait for Clk_period;
		Addr <=  "00000000010010";
		Trees_din <= x"00a400ed";
		wait for Clk_period;
		Addr <=  "00000000010011";
		Trees_din <= x"ff7500ed";
		wait for Clk_period;
		Addr <=  "00000000010100";
		Trees_din <= x"1200a004";
		wait for Clk_period;
		Addr <=  "00000000010101";
		Trees_din <= x"02e100ed";
		wait for Clk_period;
		Addr <=  "00000000010110";
		Trees_din <= x"ff9d00ed";
		wait for Clk_period;
		Addr <=  "00000000010111";
		Trees_din <= x"000c1010";
		wait for Clk_period;
		Addr <=  "00000000011000";
		Trees_din <= x"00f56608";
		wait for Clk_period;
		Addr <=  "00000000011001";
		Trees_din <= x"03fd1f04";
		wait for Clk_period;
		Addr <=  "00000000011010";
		Trees_din <= x"002700ed";
		wait for Clk_period;
		Addr <=  "00000000011011";
		Trees_din <= x"ff5b00ed";
		wait for Clk_period;
		Addr <=  "00000000011100";
		Trees_din <= x"02fcdf04";
		wait for Clk_period;
		Addr <=  "00000000011101";
		Trees_din <= x"000000ed";
		wait for Clk_period;
		Addr <=  "00000000011110";
		Trees_din <= x"029f00ed";
		wait for Clk_period;
		Addr <=  "00000000011111";
		Trees_din <= x"02ff8c04";
		wait for Clk_period;
		Addr <=  "00000000100000";
		Trees_din <= x"ff5500ed";
		wait for Clk_period;
		Addr <=  "00000000100001";
		Trees_din <= x"01f9cc04";
		wait for Clk_period;
		Addr <=  "00000000100010";
		Trees_din <= x"ff8900ed";
		wait for Clk_period;
		Addr <=  "00000000100011";
		Trees_din <= x"002700ed";
		wait for Clk_period;
		Addr <=  "00000000100100";
		Trees_din <= x"02107428";
		wait for Clk_period;
		Addr <=  "00000000100101";
		Trees_din <= x"000c1010";
		wait for Clk_period;
		Addr <=  "00000000100110";
		Trees_din <= x"0118430c";
		wait for Clk_period;
		Addr <=  "00000000100111";
		Trees_din <= x"040ac904";
		wait for Clk_period;
		Addr <=  "00000000101000";
		Trees_din <= x"042100ed";
		wait for Clk_period;
		Addr <=  "00000000101001";
		Trees_din <= x"05109304";
		wait for Clk_period;
		Addr <=  "00000000101010";
		Trees_din <= x"ff9d00ed";
		wait for Clk_period;
		Addr <=  "00000000101011";
		Trees_din <= x"028000ed";
		wait for Clk_period;
		Addr <=  "00000000101100";
		Trees_din <= x"ff8900ed";
		wait for Clk_period;
		Addr <=  "00000000101101";
		Trees_din <= x"03fcf110";
		wait for Clk_period;
		Addr <=  "00000000101110";
		Trees_din <= x"1b01d808";
		wait for Clk_period;
		Addr <=  "00000000101111";
		Trees_din <= x"08005304";
		wait for Clk_period;
		Addr <=  "00000000110000";
		Trees_din <= x"00b200ed";
		wait for Clk_period;
		Addr <=  "00000000110001";
		Trees_din <= x"028000ed";
		wait for Clk_period;
		Addr <=  "00000000110010";
		Trees_din <= x"000de204";
		wait for Clk_period;
		Addr <=  "00000000110011";
		Trees_din <= x"00b200ed";
		wait for Clk_period;
		Addr <=  "00000000110100";
		Trees_din <= x"ff9d00ed";
		wait for Clk_period;
		Addr <=  "00000000110101";
		Trees_din <= x"08005604";
		wait for Clk_period;
		Addr <=  "00000000110110";
		Trees_din <= x"ff7500ed";
		wait for Clk_period;
		Addr <=  "00000000110111";
		Trees_din <= x"002700ed";
		wait for Clk_period;
		Addr <=  "00000000111000";
		Trees_din <= x"0515e904";
		wait for Clk_period;
		Addr <=  "00000000111001";
		Trees_din <= x"ff5e00ed";
		wait for Clk_period;
		Addr <=  "00000000111010";
		Trees_din <= x"023600ed";
		wait for Clk_period;
		Addr <=  "00000000111011";
		Trees_din <= x"0509dd40";
		wait for Clk_period;
		Addr <=  "00000000111100";
		Trees_din <= x"05081c1c";
		wait for Clk_period;
		Addr <=  "00000000111101";
		Trees_din <= x"0506f70c";
		wait for Clk_period;
		Addr <=  "00000000111110";
		Trees_din <= x"20000e04";
		wait for Clk_period;
		Addr <=  "00000000111111";
		Trees_din <= x"ff5501c9";
		wait for Clk_period;
		Addr <=  "00000001000000";
		Trees_din <= x"07005504";
		wait for Clk_period;
		Addr <=  "00000001000001";
		Trees_din <= x"ff7b01c9";
		wait for Clk_period;
		Addr <=  "00000001000010";
		Trees_din <= x"003a01c9";
		wait for Clk_period;
		Addr <=  "00000001000011";
		Trees_din <= x"0d03eb08";
		wait for Clk_period;
		Addr <=  "00000001000100";
		Trees_din <= x"1304c504";
		wait for Clk_period;
		Addr <=  "00000001000101";
		Trees_din <= x"ff5901c9";
		wait for Clk_period;
		Addr <=  "00000001000110";
		Trees_din <= x"002501c9";
		wait for Clk_period;
		Addr <=  "00000001000111";
		Trees_din <= x"03fc9c04";
		wait for Clk_period;
		Addr <=  "00000001001000";
		Trees_din <= x"015c01c9";
		wait for Clk_period;
		Addr <=  "00000001001001";
		Trees_din <= x"ff9201c9";
		wait for Clk_period;
		Addr <=  "00000001001010";
		Trees_din <= x"03fb5908";
		wait for Clk_period;
		Addr <=  "00000001001011";
		Trees_din <= x"02051104";
		wait for Clk_period;
		Addr <=  "00000001001100";
		Trees_din <= x"018301c9";
		wait for Clk_period;
		Addr <=  "00000001001101";
		Trees_din <= x"ff8f01c9";
		wait for Clk_period;
		Addr <=  "00000001001110";
		Trees_din <= x"04feaa10";
		wait for Clk_period;
		Addr <=  "00000001001111";
		Trees_din <= x"0201d908";
		wait for Clk_period;
		Addr <=  "00000001010000";
		Trees_din <= x"08005704";
		wait for Clk_period;
		Addr <=  "00000001010001";
		Trees_din <= x"ff6901c9";
		wait for Clk_period;
		Addr <=  "00000001010010";
		Trees_din <= x"005601c9";
		wait for Clk_period;
		Addr <=  "00000001010011";
		Trees_din <= x"1503f004";
		wait for Clk_period;
		Addr <=  "00000001010100";
		Trees_din <= x"017b01c9";
		wait for Clk_period;
		Addr <=  "00000001010101";
		Trees_din <= x"002601c9";
		wait for Clk_period;
		Addr <=  "00000001010110";
		Trees_din <= x"0bf97704";
		wait for Clk_period;
		Addr <=  "00000001010111";
		Trees_din <= x"006501c9";
		wait for Clk_period;
		Addr <=  "00000001011000";
		Trees_din <= x"08004704";
		wait for Clk_period;
		Addr <=  "00000001011001";
		Trees_din <= x"002a01c9";
		wait for Clk_period;
		Addr <=  "00000001011010";
		Trees_din <= x"ff5b01c9";
		wait for Clk_period;
		Addr <=  "00000001011011";
		Trees_din <= x"000c631c";
		wait for Clk_period;
		Addr <=  "00000001011100";
		Trees_din <= x"0216d914";
		wait for Clk_period;
		Addr <=  "00000001011101";
		Trees_din <= x"01184310";
		wait for Clk_period;
		Addr <=  "00000001011110";
		Trees_din <= x"000b0b08";
		wait for Clk_period;
		Addr <=  "00000001011111";
		Trees_din <= x"07006004";
		wait for Clk_period;
		Addr <=  "00000001100000";
		Trees_din <= x"01ac01c9";
		wait for Clk_period;
		Addr <=  "00000001100001";
		Trees_din <= x"008d01c9";
		wait for Clk_period;
		Addr <=  "00000001100010";
		Trees_din <= x"0b022b04";
		wait for Clk_period;
		Addr <=  "00000001100011";
		Trees_din <= x"016a01c9";
		wait for Clk_period;
		Addr <=  "00000001100100";
		Trees_din <= x"003301c9";
		wait for Clk_period;
		Addr <=  "00000001100101";
		Trees_din <= x"ff7b01c9";
		wait for Clk_period;
		Addr <=  "00000001100110";
		Trees_din <= x"1900a704";
		wait for Clk_period;
		Addr <=  "00000001100111";
		Trees_din <= x"ff6701c9";
		wait for Clk_period;
		Addr <=  "00000001101000";
		Trees_din <= x"002f01c9";
		wait for Clk_period;
		Addr <=  "00000001101001";
		Trees_din <= x"03fcc70c";
		wait for Clk_period;
		Addr <=  "00000001101010";
		Trees_din <= x"000e8708";
		wait for Clk_period;
		Addr <=  "00000001101011";
		Trees_din <= x"1000de04";
		wait for Clk_period;
		Addr <=  "00000001101100";
		Trees_din <= x"01b301c9";
		wait for Clk_period;
		Addr <=  "00000001101101";
		Trees_din <= x"007c01c9";
		wait for Clk_period;
		Addr <=  "00000001101110";
		Trees_din <= x"ff9a01c9";
		wait for Clk_period;
		Addr <=  "00000001101111";
		Trees_din <= x"07005b04";
		wait for Clk_period;
		Addr <=  "00000001110000";
		Trees_din <= x"ff6501c9";
		wait for Clk_period;
		Addr <=  "00000001110001";
		Trees_din <= x"003c01c9";
		wait for Clk_period;
		Addr <=  "00000001110010";
		Trees_din <= x"0509dd34";
		wait for Clk_period;
		Addr <=  "00000001110011";
		Trees_din <= x"05081c1c";
		wait for Clk_period;
		Addr <=  "00000001110100";
		Trees_din <= x"0506f70c";
		wait for Clk_period;
		Addr <=  "00000001110101";
		Trees_din <= x"20000e04";
		wait for Clk_period;
		Addr <=  "00000001110110";
		Trees_din <= x"ff590275";
		wait for Clk_period;
		Addr <=  "00000001110111";
		Trees_din <= x"13fb1304";
		wait for Clk_period;
		Addr <=  "00000001111000";
		Trees_din <= x"003b0275";
		wait for Clk_period;
		Addr <=  "00000001111001";
		Trees_din <= x"ff840275";
		wait for Clk_period;
		Addr <=  "00000001111010";
		Trees_din <= x"0d03eb08";
		wait for Clk_period;
		Addr <=  "00000001111011";
		Trees_din <= x"04fd7604";
		wait for Clk_period;
		Addr <=  "00000001111100";
		Trees_din <= x"00280275";
		wait for Clk_period;
		Addr <=  "00000001111101";
		Trees_din <= x"ff5f0275";
		wait for Clk_period;
		Addr <=  "00000001111110";
		Trees_din <= x"0f022704";
		wait for Clk_period;
		Addr <=  "00000001111111";
		Trees_din <= x"ff9a0275";
		wait for Clk_period;
		Addr <=  "00000010000000";
		Trees_din <= x"010e0275";
		wait for Clk_period;
		Addr <=  "00000010000001";
		Trees_din <= x"000e4210";
		wait for Clk_period;
		Addr <=  "00000010000010";
		Trees_din <= x"00f56604";
		wait for Clk_period;
		Addr <=  "00000010000011";
		Trees_din <= x"ff660275";
		wait for Clk_period;
		Addr <=  "00000010000100";
		Trees_din <= x"0ef8ee04";
		wait for Clk_period;
		Addr <=  "00000010000101";
		Trees_din <= x"ff8e0275";
		wait for Clk_period;
		Addr <=  "00000010000110";
		Trees_din <= x"02fced04";
		wait for Clk_period;
		Addr <=  "00000010000111";
		Trees_din <= x"ffe80275";
		wait for Clk_period;
		Addr <=  "00000010001000";
		Trees_din <= x"01480275";
		wait for Clk_period;
		Addr <=  "00000010001001";
		Trees_din <= x"1a005704";
		wait for Clk_period;
		Addr <=  "00000010001010";
		Trees_din <= x"ff620275";
		wait for Clk_period;
		Addr <=  "00000010001011";
		Trees_din <= x"00240275";
		wait for Clk_period;
		Addr <=  "00000010001100";
		Trees_din <= x"0216d91c";
		wait for Clk_period;
		Addr <=  "00000010001101";
		Trees_din <= x"000d8d10";
		wait for Clk_period;
		Addr <=  "00000010001110";
		Trees_din <= x"0118430c";
		wait for Clk_period;
		Addr <=  "00000010001111";
		Trees_din <= x"000b0b04";
		wait for Clk_period;
		Addr <=  "00000010010000";
		Trees_din <= x"01310275";
		wait for Clk_period;
		Addr <=  "00000010010001";
		Trees_din <= x"03fcf104";
		wait for Clk_period;
		Addr <=  "00000010010010";
		Trees_din <= x"011a0275";
		wait for Clk_period;
		Addr <=  "00000010010011";
		Trees_din <= x"000b0275";
		wait for Clk_period;
		Addr <=  "00000010010100";
		Trees_din <= x"ff840275";
		wait for Clk_period;
		Addr <=  "00000010010101";
		Trees_din <= x"03fc9208";
		wait for Clk_period;
		Addr <=  "00000010010110";
		Trees_din <= x"1101b504";
		wait for Clk_period;
		Addr <=  "00000010010111";
		Trees_din <= x"ffa60275";
		wait for Clk_period;
		Addr <=  "00000010011000";
		Trees_din <= x"00fd0275";
		wait for Clk_period;
		Addr <=  "00000010011001";
		Trees_din <= x"ff6e0275";
		wait for Clk_period;
		Addr <=  "00000010011010";
		Trees_din <= x"09059704";
		wait for Clk_period;
		Addr <=  "00000010011011";
		Trees_din <= x"ff6e0275";
		wait for Clk_period;
		Addr <=  "00000010011100";
		Trees_din <= x"003b0275";
		wait for Clk_period;
		Addr <=  "00000010011101";
		Trees_din <= x"0509dd48";
		wait for Clk_period;
		Addr <=  "00000010011110";
		Trees_din <= x"05081c20";
		wait for Clk_period;
		Addr <=  "00000010011111";
		Trees_din <= x"0506f70c";
		wait for Clk_period;
		Addr <=  "00000010100000";
		Trees_din <= x"20000e04";
		wait for Clk_period;
		Addr <=  "00000010100001";
		Trees_din <= x"ff5d0341";
		wait for Clk_period;
		Addr <=  "00000010100010";
		Trees_din <= x"03fe1f04";
		wait for Clk_period;
		Addr <=  "00000010100011";
		Trees_din <= x"003e0341";
		wait for Clk_period;
		Addr <=  "00000010100100";
		Trees_din <= x"ff8c0341";
		wait for Clk_period;
		Addr <=  "00000010100101";
		Trees_din <= x"03fbcb0c";
		wait for Clk_period;
		Addr <=  "00000010100110";
		Trees_din <= x"17004404";
		wait for Clk_period;
		Addr <=  "00000010100111";
		Trees_din <= x"ffa00341";
		wait for Clk_period;
		Addr <=  "00000010101000";
		Trees_din <= x"0eff8804";
		wait for Clk_period;
		Addr <=  "00000010101001";
		Trees_din <= x"01240341";
		wait for Clk_period;
		Addr <=  "00000010101010";
		Trees_din <= x"00290341";
		wait for Clk_period;
		Addr <=  "00000010101011";
		Trees_din <= x"17005004";
		wait for Clk_period;
		Addr <=  "00000010101100";
		Trees_din <= x"ff630341";
		wait for Clk_period;
		Addr <=  "00000010101101";
		Trees_din <= x"001b0341";
		wait for Clk_period;
		Addr <=  "00000010101110";
		Trees_din <= x"03fc6b10";
		wait for Clk_period;
		Addr <=  "00000010101111";
		Trees_din <= x"14034c0c";
		wait for Clk_period;
		Addr <=  "00000010110000";
		Trees_din <= x"10fe2904";
		wait for Clk_period;
		Addr <=  "00000010110001";
		Trees_din <= x"ffa30341";
		wait for Clk_period;
		Addr <=  "00000010110010";
		Trees_din <= x"17003e04";
		wait for Clk_period;
		Addr <=  "00000010110011";
		Trees_din <= x"002c0341";
		wait for Clk_period;
		Addr <=  "00000010110100";
		Trees_din <= x"013d0341";
		wait for Clk_period;
		Addr <=  "00000010110101";
		Trees_din <= x"ff890341";
		wait for Clk_period;
		Addr <=  "00000010110110";
		Trees_din <= x"04fe610c";
		wait for Clk_period;
		Addr <=  "00000010110111";
		Trees_din <= x"000e0608";
		wait for Clk_period;
		Addr <=  "00000010111000";
		Trees_din <= x"19009c04";
		wait for Clk_period;
		Addr <=  "00000010111001";
		Trees_din <= x"fffc0341";
		wait for Clk_period;
		Addr <=  "00000010111010";
		Trees_din <= x"00ff0341";
		wait for Clk_period;
		Addr <=  "00000010111011";
		Trees_din <= x"ff960341";
		wait for Clk_period;
		Addr <=  "00000010111100";
		Trees_din <= x"20000008";
		wait for Clk_period;
		Addr <=  "00000010111101";
		Trees_din <= x"0ffc5f04";
		wait for Clk_period;
		Addr <=  "00000010111110";
		Trees_din <= x"00250341";
		wait for Clk_period;
		Addr <=  "00000010111111";
		Trees_din <= x"ff640341";
		wait for Clk_period;
		Addr <=  "00000011000000";
		Trees_din <= x"00550341";
		wait for Clk_period;
		Addr <=  "00000011000001";
		Trees_din <= x"02107418";
		wait for Clk_period;
		Addr <=  "00000011000010";
		Trees_din <= x"000de210";
		wait for Clk_period;
		Addr <=  "00000011000011";
		Trees_din <= x"0118430c";
		wait for Clk_period;
		Addr <=  "00000011000100";
		Trees_din <= x"000b0b04";
		wait for Clk_period;
		Addr <=  "00000011000101";
		Trees_din <= x"00f80341";
		wait for Clk_period;
		Addr <=  "00000011000110";
		Trees_din <= x"03fcf104";
		wait for Clk_period;
		Addr <=  "00000011000111";
		Trees_din <= x"00e60341";
		wait for Clk_period;
		Addr <=  "00000011001000";
		Trees_din <= x"fff50341";
		wait for Clk_period;
		Addr <=  "00000011001001";
		Trees_din <= x"ffa50341";
		wait for Clk_period;
		Addr <=  "00000011001010";
		Trees_din <= x"08005904";
		wait for Clk_period;
		Addr <=  "00000011001011";
		Trees_din <= x"ff740341";
		wait for Clk_period;
		Addr <=  "00000011001100";
		Trees_din <= x"00750341";
		wait for Clk_period;
		Addr <=  "00000011001101";
		Trees_din <= x"0515e904";
		wait for Clk_period;
		Addr <=  "00000011001110";
		Trees_din <= x"ff6b0341";
		wait for Clk_period;
		Addr <=  "00000011001111";
		Trees_din <= x"00e40341";
		wait for Clk_period;
		Addr <=  "00000011010000";
		Trees_din <= x"0509dd40";
		wait for Clk_period;
		Addr <=  "00000011010001";
		Trees_din <= x"05072414";
		wait for Clk_period;
		Addr <=  "00000011010010";
		Trees_din <= x"20000e0c";
		wait for Clk_period;
		Addr <=  "00000011010011";
		Trees_din <= x"0506f704";
		wait for Clk_period;
		Addr <=  "00000011010100";
		Trees_din <= x"ff600425";
		wait for Clk_period;
		Addr <=  "00000011010101";
		Trees_din <= x"11003904";
		wait for Clk_period;
		Addr <=  "00000011010110";
		Trees_din <= x"002b0425";
		wait for Clk_period;
		Addr <=  "00000011010111";
		Trees_din <= x"ff850425";
		wait for Clk_period;
		Addr <=  "00000011011000";
		Trees_din <= x"0200c104";
		wait for Clk_period;
		Addr <=  "00000011011001";
		Trees_din <= x"ff950425";
		wait for Clk_period;
		Addr <=  "00000011011010";
		Trees_din <= x"00390425";
		wait for Clk_period;
		Addr <=  "00000011011011";
		Trees_din <= x"03fbd814";
		wait for Clk_period;
		Addr <=  "00000011011100";
		Trees_din <= x"1c003208";
		wait for Clk_period;
		Addr <=  "00000011011101";
		Trees_din <= x"1d00e004";
		wait for Clk_period;
		Addr <=  "00000011011110";
		Trees_din <= x"ff8a0425";
		wait for Clk_period;
		Addr <=  "00000011011111";
		Trees_din <= x"00280425";
		wait for Clk_period;
		Addr <=  "00000011100000";
		Trees_din <= x"0a006404";
		wait for Clk_period;
		Addr <=  "00000011100001";
		Trees_din <= x"000a0425";
		wait for Clk_period;
		Addr <=  "00000011100010";
		Trees_din <= x"17004404";
		wait for Clk_period;
		Addr <=  "00000011100011";
		Trees_din <= x"00570425";
		wait for Clk_period;
		Addr <=  "00000011100100";
		Trees_din <= x"014d0425";
		wait for Clk_period;
		Addr <=  "00000011100101";
		Trees_din <= x"04fe610c";
		wait for Clk_period;
		Addr <=  "00000011100110";
		Trees_din <= x"000e0608";
		wait for Clk_period;
		Addr <=  "00000011100111";
		Trees_din <= x"01fa6304";
		wait for Clk_period;
		Addr <=  "00000011101000";
		Trees_din <= x"ffcc0425";
		wait for Clk_period;
		Addr <=  "00000011101001";
		Trees_din <= x"00eb0425";
		wait for Clk_period;
		Addr <=  "00000011101010";
		Trees_din <= x"ff850425";
		wait for Clk_period;
		Addr <=  "00000011101011";
		Trees_din <= x"18005308";
		wait for Clk_period;
		Addr <=  "00000011101100";
		Trees_din <= x"20000004";
		wait for Clk_period;
		Addr <=  "00000011101101";
		Trees_din <= x"ff640425";
		wait for Clk_period;
		Addr <=  "00000011101110";
		Trees_din <= x"00330425";
		wait for Clk_period;
		Addr <=  "00000011101111";
		Trees_din <= x"00820425";
		wait for Clk_period;
		Addr <=  "00000011110000";
		Trees_din <= x"050d5a20";
		wait for Clk_period;
		Addr <=  "00000011110001";
		Trees_din <= x"00ddf604";
		wait for Clk_period;
		Addr <=  "00000011110010";
		Trees_din <= x"ff6c0425";
		wait for Clk_period;
		Addr <=  "00000011110011";
		Trees_din <= x"000c100c";
		wait for Clk_period;
		Addr <=  "00000011110100";
		Trees_din <= x"02faea04";
		wait for Clk_period;
		Addr <=  "00000011110101";
		Trees_din <= x"ff700425";
		wait for Clk_period;
		Addr <=  "00000011110110";
		Trees_din <= x"020c5e04";
		wait for Clk_period;
		Addr <=  "00000011110111";
		Trees_din <= x"00cc0425";
		wait for Clk_period;
		Addr <=  "00000011111000";
		Trees_din <= x"ff8b0425";
		wait for Clk_period;
		Addr <=  "00000011111001";
		Trees_din <= x"08005808";
		wait for Clk_period;
		Addr <=  "00000011111010";
		Trees_din <= x"1c002504";
		wait for Clk_period;
		Addr <=  "00000011111011";
		Trees_din <= x"00330425";
		wait for Clk_period;
		Addr <=  "00000011111100";
		Trees_din <= x"ff690425";
		wait for Clk_period;
		Addr <=  "00000011111101";
		Trees_din <= x"08005904";
		wait for Clk_period;
		Addr <=  "00000011111110";
		Trees_din <= x"00fb0425";
		wait for Clk_period;
		Addr <=  "00000011111111";
		Trees_din <= x"000c0425";
		wait for Clk_period;
		Addr <=  "00000100000000";
		Trees_din <= x"021b0610";
		wait for Clk_period;
		Addr <=  "00000100000001";
		Trees_din <= x"0118430c";
		wait for Clk_period;
		Addr <=  "00000100000010";
		Trees_din <= x"000de208";
		wait for Clk_period;
		Addr <=  "00000100000011";
		Trees_din <= x"07006004";
		wait for Clk_period;
		Addr <=  "00000100000100";
		Trees_din <= x"00db0425";
		wait for Clk_period;
		Addr <=  "00000100000101";
		Trees_din <= x"00380425";
		wait for Clk_period;
		Addr <=  "00000100000110";
		Trees_din <= x"00250425";
		wait for Clk_period;
		Addr <=  "00000100000111";
		Trees_din <= x"00040425";
		wait for Clk_period;
		Addr <=  "00000100001000";
		Trees_din <= x"ff950425";
		wait for Clk_period;
		Addr <=  "00000100001001";
		Trees_din <= x"05085530";
		wait for Clk_period;
		Addr <=  "00000100001010";
		Trees_din <= x"0506f718";
		wait for Clk_period;
		Addr <=  "00000100001011";
		Trees_din <= x"20000e10";
		wait for Clk_period;
		Addr <=  "00000100001100";
		Trees_din <= x"10040c04";
		wait for Clk_period;
		Addr <=  "00000100001101";
		Trees_din <= x"ff6104f9";
		wait for Clk_period;
		Addr <=  "00000100001110";
		Trees_din <= x"05039504";
		wait for Clk_period;
		Addr <=  "00000100001111";
		Trees_din <= x"ff6a04f9";
		wait for Clk_period;
		Addr <=  "00000100010000";
		Trees_din <= x"0a02ce04";
		wait for Clk_period;
		Addr <=  "00000100010001";
		Trees_din <= x"ff9904f9";
		wait for Clk_period;
		Addr <=  "00000100010010";
		Trees_din <= x"00de04f9";
		wait for Clk_period;
		Addr <=  "00000100010011";
		Trees_din <= x"08005504";
		wait for Clk_period;
		Addr <=  "00000100010100";
		Trees_din <= x"ff9d04f9";
		wait for Clk_period;
		Addr <=  "00000100010101";
		Trees_din <= x"003904f9";
		wait for Clk_period;
		Addr <=  "00000100010110";
		Trees_din <= x"03fbcb0c";
		wait for Clk_period;
		Addr <=  "00000100010111";
		Trees_din <= x"0d023004";
		wait for Clk_period;
		Addr <=  "00000100011000";
		Trees_din <= x"ffa004f9";
		wait for Clk_period;
		Addr <=  "00000100011001";
		Trees_din <= x"17004404";
		wait for Clk_period;
		Addr <=  "00000100011010";
		Trees_din <= x"001004f9";
		wait for Clk_period;
		Addr <=  "00000100011011";
		Trees_din <= x"00e004f9";
		wait for Clk_period;
		Addr <=  "00000100011100";
		Trees_din <= x"04fe2208";
		wait for Clk_period;
		Addr <=  "00000100011101";
		Trees_din <= x"15f97c04";
		wait for Clk_period;
		Addr <=  "00000100011110";
		Trees_din <= x"006604f9";
		wait for Clk_period;
		Addr <=  "00000100011111";
		Trees_din <= x"ff9a04f9";
		wait for Clk_period;
		Addr <=  "00000100100000";
		Trees_din <= x"ff6b04f9";
		wait for Clk_period;
		Addr <=  "00000100100001";
		Trees_din <= x"050d5a28";
		wait for Clk_period;
		Addr <=  "00000100100010";
		Trees_din <= x"03fcf114";
		wait for Clk_period;
		Addr <=  "00000100100011";
		Trees_din <= x"020c5e10";
		wait for Clk_period;
		Addr <=  "00000100100100";
		Trees_din <= x"000e6e08";
		wait for Clk_period;
		Addr <=  "00000100100101";
		Trees_din <= x"0a000504";
		wait for Clk_period;
		Addr <=  "00000100100110";
		Trees_din <= x"ffce04f9";
		wait for Clk_period;
		Addr <=  "00000100100111";
		Trees_din <= x"00c804f9";
		wait for Clk_period;
		Addr <=  "00000100101000";
		Trees_din <= x"1b038604";
		wait for Clk_period;
		Addr <=  "00000100101001";
		Trees_din <= x"ff8c04f9";
		wait for Clk_period;
		Addr <=  "00000100101010";
		Trees_din <= x"003304f9";
		wait for Clk_period;
		Addr <=  "00000100101011";
		Trees_din <= x"ff8204f9";
		wait for Clk_period;
		Addr <=  "00000100101100";
		Trees_din <= x"00ec0004";
		wait for Clk_period;
		Addr <=  "00000100101101";
		Trees_din <= x"ff6704f9";
		wait for Clk_period;
		Addr <=  "00000100101110";
		Trees_din <= x"0008f408";
		wait for Clk_period;
		Addr <=  "00000100101111";
		Trees_din <= x"00f56604";
		wait for Clk_period;
		Addr <=  "00000100110000";
		Trees_din <= x"000104f9";
		wait for Clk_period;
		Addr <=  "00000100110001";
		Trees_din <= x"00b304f9";
		wait for Clk_period;
		Addr <=  "00000100110010";
		Trees_din <= x"09f96b04";
		wait for Clk_period;
		Addr <=  "00000100110011";
		Trees_din <= x"00b404f9";
		wait for Clk_period;
		Addr <=  "00000100110100";
		Trees_din <= x"ff8404f9";
		wait for Clk_period;
		Addr <=  "00000100110101";
		Trees_din <= x"021b0610";
		wait for Clk_period;
		Addr <=  "00000100110110";
		Trees_din <= x"0118430c";
		wait for Clk_period;
		Addr <=  "00000100110111";
		Trees_din <= x"07006008";
		wait for Clk_period;
		Addr <=  "00000100111000";
		Trees_din <= x"040db704";
		wait for Clk_period;
		Addr <=  "00000100111001";
		Trees_din <= x"00c604f9";
		wait for Clk_period;
		Addr <=  "00000100111010";
		Trees_din <= x"003704f9";
		wait for Clk_period;
		Addr <=  "00000100111011";
		Trees_din <= x"003004f9";
		wait for Clk_period;
		Addr <=  "00000100111100";
		Trees_din <= x"000a04f9";
		wait for Clk_period;
		Addr <=  "00000100111101";
		Trees_din <= x"ff9c04f9";
		wait for Clk_period;
		Addr <=  "00000100111110";
		Trees_din <= x"0508552c";
		wait for Clk_period;
		Addr <=  "00000100111111";
		Trees_din <= x"0506f718";
		wait for Clk_period;
		Addr <=  "00000101000000";
		Trees_din <= x"20000e10";
		wait for Clk_period;
		Addr <=  "00000101000001";
		Trees_din <= x"10040c04";
		wait for Clk_period;
		Addr <=  "00000101000010";
		Trees_din <= x"ff6305c5";
		wait for Clk_period;
		Addr <=  "00000101000011";
		Trees_din <= x"05039504";
		wait for Clk_period;
		Addr <=  "00000101000100";
		Trees_din <= x"ff6d05c5";
		wait for Clk_period;
		Addr <=  "00000101000101";
		Trees_din <= x"05044004";
		wait for Clk_period;
		Addr <=  "00000101000110";
		Trees_din <= x"00d705c5";
		wait for Clk_period;
		Addr <=  "00000101000111";
		Trees_din <= x"ff9e05c5";
		wait for Clk_period;
		Addr <=  "00000101001000";
		Trees_din <= x"17004304";
		wait for Clk_period;
		Addr <=  "00000101001001";
		Trees_din <= x"ffa605c5";
		wait for Clk_period;
		Addr <=  "00000101001010";
		Trees_din <= x"003405c5";
		wait for Clk_period;
		Addr <=  "00000101001011";
		Trees_din <= x"1400520c";
		wait for Clk_period;
		Addr <=  "00000101001100";
		Trees_din <= x"03fc9c08";
		wait for Clk_period;
		Addr <=  "00000101001101";
		Trees_din <= x"04fe5004";
		wait for Clk_period;
		Addr <=  "00000101001110";
		Trees_din <= x"00c105c5";
		wait for Clk_period;
		Addr <=  "00000101001111";
		Trees_din <= x"000e05c5";
		wait for Clk_period;
		Addr <=  "00000101010000";
		Trees_din <= x"ff9505c5";
		wait for Clk_period;
		Addr <=  "00000101010001";
		Trees_din <= x"0a000704";
		wait for Clk_period;
		Addr <=  "00000101010010";
		Trees_din <= x"ffeb05c5";
		wait for Clk_period;
		Addr <=  "00000101010011";
		Trees_din <= x"ff6f05c5";
		wait for Clk_period;
		Addr <=  "00000101010100";
		Trees_din <= x"050d5a24";
		wait for Clk_period;
		Addr <=  "00000101010101";
		Trees_din <= x"00f4590c";
		wait for Clk_period;
		Addr <=  "00000101010110";
		Trees_din <= x"03fd1f08";
		wait for Clk_period;
		Addr <=  "00000101010111";
		Trees_din <= x"19008c04";
		wait for Clk_period;
		Addr <=  "00000101011000";
		Trees_din <= x"006e05c5";
		wait for Clk_period;
		Addr <=  "00000101011001";
		Trees_din <= x"ffa105c5";
		wait for Clk_period;
		Addr <=  "00000101011010";
		Trees_din <= x"ff6c05c5";
		wait for Clk_period;
		Addr <=  "00000101011011";
		Trees_din <= x"000e6e10";
		wait for Clk_period;
		Addr <=  "00000101011100";
		Trees_din <= x"0ef8f708";
		wait for Clk_period;
		Addr <=  "00000101011101";
		Trees_din <= x"14022804";
		wait for Clk_period;
		Addr <=  "00000101011110";
		Trees_din <= x"005e05c5";
		wait for Clk_period;
		Addr <=  "00000101011111";
		Trees_din <= x"ff8905c5";
		wait for Clk_period;
		Addr <=  "00000101100000";
		Trees_din <= x"02fa1e04";
		wait for Clk_period;
		Addr <=  "00000101100001";
		Trees_din <= x"ff9f05c5";
		wait for Clk_period;
		Addr <=  "00000101100010";
		Trees_din <= x"009b05c5";
		wait for Clk_period;
		Addr <=  "00000101100011";
		Trees_din <= x"1e008704";
		wait for Clk_period;
		Addr <=  "00000101100100";
		Trees_din <= x"ff7405c5";
		wait for Clk_period;
		Addr <=  "00000101100101";
		Trees_din <= x"002f05c5";
		wait for Clk_period;
		Addr <=  "00000101100110";
		Trees_din <= x"021b0614";
		wait for Clk_period;
		Addr <=  "00000101100111";
		Trees_din <= x"01184310";
		wait for Clk_period;
		Addr <=  "00000101101000";
		Trees_din <= x"000b0b08";
		wait for Clk_period;
		Addr <=  "00000101101001";
		Trees_din <= x"07006004";
		wait for Clk_period;
		Addr <=  "00000101101010";
		Trees_din <= x"00b905c5";
		wait for Clk_period;
		Addr <=  "00000101101011";
		Trees_din <= x"002b05c5";
		wait for Clk_period;
		Addr <=  "00000101101100";
		Trees_din <= x"03fcc704";
		wait for Clk_period;
		Addr <=  "00000101101101";
		Trees_din <= x"00a505c5";
		wait for Clk_period;
		Addr <=  "00000101101110";
		Trees_din <= x"ffe205c5";
		wait for Clk_period;
		Addr <=  "00000101101111";
		Trees_din <= x"000d05c5";
		wait for Clk_period;
		Addr <=  "00000101110000";
		Trees_din <= x"ffa405c5";
		wait for Clk_period;
		Addr <=  "00000101110001";
		Trees_din <= x"05085528";
		wait for Clk_period;
		Addr <=  "00000101110010";
		Trees_din <= x"0506f714";
		wait for Clk_period;
		Addr <=  "00000101110011";
		Trees_din <= x"20000e10";
		wait for Clk_period;
		Addr <=  "00000101110100";
		Trees_din <= x"10040c04";
		wait for Clk_period;
		Addr <=  "00000101110101";
		Trees_din <= x"ff640679";
		wait for Clk_period;
		Addr <=  "00000101110110";
		Trees_din <= x"05039504";
		wait for Clk_period;
		Addr <=  "00000101110111";
		Trees_din <= x"ff720679";
		wait for Clk_period;
		Addr <=  "00000101111000";
		Trees_din <= x"06fe5004";
		wait for Clk_period;
		Addr <=  "00000101111001";
		Trees_din <= x"ffa20679";
		wait for Clk_period;
		Addr <=  "00000101111010";
		Trees_din <= x"00d30679";
		wait for Clk_period;
		Addr <=  "00000101111011";
		Trees_din <= x"ffea0679";
		wait for Clk_period;
		Addr <=  "00000101111100";
		Trees_din <= x"1400520c";
		wait for Clk_period;
		Addr <=  "00000101111101";
		Trees_din <= x"03fc9c08";
		wait for Clk_period;
		Addr <=  "00000101111110";
		Trees_din <= x"1f028804";
		wait for Clk_period;
		Addr <=  "00000101111111";
		Trees_din <= x"00030679";
		wait for Clk_period;
		Addr <=  "00000110000000";
		Trees_din <= x"00b00679";
		wait for Clk_period;
		Addr <=  "00000110000001";
		Trees_din <= x"ff9e0679";
		wait for Clk_period;
		Addr <=  "00000110000010";
		Trees_din <= x"06fb9204";
		wait for Clk_period;
		Addr <=  "00000110000011";
		Trees_din <= x"fff20679";
		wait for Clk_period;
		Addr <=  "00000110000100";
		Trees_din <= x"ff740679";
		wait for Clk_period;
		Addr <=  "00000110000101";
		Trees_din <= x"050d5a1c";
		wait for Clk_period;
		Addr <=  "00000110000110";
		Trees_din <= x"020c5e18";
		wait for Clk_period;
		Addr <=  "00000110000111";
		Trees_din <= x"000e6e10";
		wait for Clk_period;
		Addr <=  "00000110001000";
		Trees_din <= x"03fd6008";
		wait for Clk_period;
		Addr <=  "00000110001001";
		Trees_din <= x"01fa0c04";
		wait for Clk_period;
		Addr <=  "00000110001010";
		Trees_din <= x"000d0679";
		wait for Clk_period;
		Addr <=  "00000110001011";
		Trees_din <= x"00a10679";
		wait for Clk_period;
		Addr <=  "00000110001100";
		Trees_din <= x"04002a04";
		wait for Clk_period;
		Addr <=  "00000110001101";
		Trees_din <= x"00400679";
		wait for Clk_period;
		Addr <=  "00000110001110";
		Trees_din <= x"ff980679";
		wait for Clk_period;
		Addr <=  "00000110001111";
		Trees_din <= x"0c001a04";
		wait for Clk_period;
		Addr <=  "00000110010000";
		Trees_din <= x"002c0679";
		wait for Clk_period;
		Addr <=  "00000110010001";
		Trees_din <= x"ff790679";
		wait for Clk_period;
		Addr <=  "00000110010010";
		Trees_din <= x"ff760679";
		wait for Clk_period;
		Addr <=  "00000110010011";
		Trees_din <= x"021b0614";
		wait for Clk_period;
		Addr <=  "00000110010100";
		Trees_din <= x"01184310";
		wait for Clk_period;
		Addr <=  "00000110010101";
		Trees_din <= x"000b0b08";
		wait for Clk_period;
		Addr <=  "00000110010110";
		Trees_din <= x"040db704";
		wait for Clk_period;
		Addr <=  "00000110010111";
		Trees_din <= x"00b00679";
		wait for Clk_period;
		Addr <=  "00000110011000";
		Trees_din <= x"001c0679";
		wait for Clk_period;
		Addr <=  "00000110011001";
		Trees_din <= x"1403ba04";
		wait for Clk_period;
		Addr <=  "00000110011010";
		Trees_din <= x"008a0679";
		wait for Clk_period;
		Addr <=  "00000110011011";
		Trees_din <= x"ffb10679";
		wait for Clk_period;
		Addr <=  "00000110011100";
		Trees_din <= x"000e0679";
		wait for Clk_period;
		Addr <=  "00000110011101";
		Trees_din <= x"ffab0679";
		wait for Clk_period;
		Addr <=  "00000110011110";
		Trees_din <= x"05085528";
		wait for Clk_period;
		Addr <=  "00000110011111";
		Trees_din <= x"0506f714";
		wait for Clk_period;
		Addr <=  "00000110100000";
		Trees_din <= x"20000e10";
		wait for Clk_period;
		Addr <=  "00000110100001";
		Trees_din <= x"10040c04";
		wait for Clk_period;
		Addr <=  "00000110100010";
		Trees_din <= x"ff66073d";
		wait for Clk_period;
		Addr <=  "00000110100011";
		Trees_din <= x"05039504";
		wait for Clk_period;
		Addr <=  "00000110100100";
		Trees_din <= x"ff76073d";
		wait for Clk_period;
		Addr <=  "00000110100101";
		Trees_din <= x"06fe7904";
		wait for Clk_period;
		Addr <=  "00000110100110";
		Trees_din <= x"ffa9073d";
		wait for Clk_period;
		Addr <=  "00000110100111";
		Trees_din <= x"00bc073d";
		wait for Clk_period;
		Addr <=  "00000110101000";
		Trees_din <= x"fff1073d";
		wait for Clk_period;
		Addr <=  "00000110101001";
		Trees_din <= x"04fe500c";
		wait for Clk_period;
		Addr <=  "00000110101010";
		Trees_din <= x"01fa8604";
		wait for Clk_period;
		Addr <=  "00000110101011";
		Trees_din <= x"ffa9073d";
		wait for Clk_period;
		Addr <=  "00000110101100";
		Trees_din <= x"12008404";
		wait for Clk_period;
		Addr <=  "00000110101101";
		Trees_din <= x"00b3073d";
		wait for Clk_period;
		Addr <=  "00000110101110";
		Trees_din <= x"0015073d";
		wait for Clk_period;
		Addr <=  "00000110101111";
		Trees_din <= x"07005b04";
		wait for Clk_period;
		Addr <=  "00000110110000";
		Trees_din <= x"ff78073d";
		wait for Clk_period;
		Addr <=  "00000110110001";
		Trees_din <= x"0005073d";
		wait for Clk_period;
		Addr <=  "00000110110010";
		Trees_din <= x"050d5a20";
		wait for Clk_period;
		Addr <=  "00000110110011";
		Trees_din <= x"00f45908";
		wait for Clk_period;
		Addr <=  "00000110110100";
		Trees_din <= x"03fd1f04";
		wait for Clk_period;
		Addr <=  "00000110110101";
		Trees_din <= x"0004073d";
		wait for Clk_period;
		Addr <=  "00000110110110";
		Trees_din <= x"ff7a073d";
		wait for Clk_period;
		Addr <=  "00000110110111";
		Trees_din <= x"000e6e10";
		wait for Clk_period;
		Addr <=  "00000110111000";
		Trees_din <= x"08005208";
		wait for Clk_period;
		Addr <=  "00000110111001";
		Trees_din <= x"0007ff04";
		wait for Clk_period;
		Addr <=  "00000110111010";
		Trees_din <= x"007a073d";
		wait for Clk_period;
		Addr <=  "00000110111011";
		Trees_din <= x"ffbc073d";
		wait for Clk_period;
		Addr <=  "00000110111100";
		Trees_din <= x"06fa6a04";
		wait for Clk_period;
		Addr <=  "00000110111101";
		Trees_din <= x"ffac073d";
		wait for Clk_period;
		Addr <=  "00000110111110";
		Trees_din <= x"0092073d";
		wait for Clk_period;
		Addr <=  "00000110111111";
		Trees_din <= x"18004a04";
		wait for Clk_period;
		Addr <=  "00000111000000";
		Trees_din <= x"ff81073d";
		wait for Clk_period;
		Addr <=  "00000111000001";
		Trees_din <= x"0022073d";
		wait for Clk_period;
		Addr <=  "00000111000010";
		Trees_din <= x"01184318";
		wait for Clk_period;
		Addr <=  "00000111000011";
		Trees_din <= x"000b0b0c";
		wait for Clk_period;
		Addr <=  "00000111000100";
		Trees_din <= x"040db708";
		wait for Clk_period;
		Addr <=  "00000111000101";
		Trees_din <= x"07006004";
		wait for Clk_period;
		Addr <=  "00000111000110";
		Trees_din <= x"00aa073d";
		wait for Clk_period;
		Addr <=  "00000111000111";
		Trees_din <= x"0015073d";
		wait for Clk_period;
		Addr <=  "00000111001000";
		Trees_din <= x"000b073d";
		wait for Clk_period;
		Addr <=  "00000111001001";
		Trees_din <= x"06fc2004";
		wait for Clk_period;
		Addr <=  "00000111001010";
		Trees_din <= x"00a2073d";
		wait for Clk_period;
		Addr <=  "00000111001011";
		Trees_din <= x"03fcc704";
		wait for Clk_period;
		Addr <=  "00000111001100";
		Trees_din <= x"004d073d";
		wait for Clk_period;
		Addr <=  "00000111001101";
		Trees_din <= x"ff83073d";
		wait for Clk_period;
		Addr <=  "00000111001110";
		Trees_din <= x"ffec073d";
		wait for Clk_period;
		Addr <=  "00000111001111";
		Trees_din <= x"05085530";
		wait for Clk_period;
		Addr <=  "00000111010000";
		Trees_din <= x"0506f71c";
		wait for Clk_period;
		Addr <=  "00000111010001";
		Trees_din <= x"21008518";
		wait for Clk_period;
		Addr <=  "00000111010010";
		Trees_din <= x"10040c0c";
		wait for Clk_period;
		Addr <=  "00000111010011";
		Trees_din <= x"15f8e908";
		wait for Clk_period;
		Addr <=  "00000111010100";
		Trees_din <= x"01fffd04";
		wait for Clk_period;
		Addr <=  "00000111010101";
		Trees_din <= x"ff7e0801";
		wait for Clk_period;
		Addr <=  "00000111010110";
		Trees_din <= x"00470801";
		wait for Clk_period;
		Addr <=  "00000111010111";
		Trees_din <= x"ff650801";
		wait for Clk_period;
		Addr <=  "00000111011000";
		Trees_din <= x"05039504";
		wait for Clk_period;
		Addr <=  "00000111011001";
		Trees_din <= x"ff7c0801";
		wait for Clk_period;
		Addr <=  "00000111011010";
		Trees_din <= x"0a02dd04";
		wait for Clk_period;
		Addr <=  "00000111011011";
		Trees_din <= x"ffb00801";
		wait for Clk_period;
		Addr <=  "00000111011100";
		Trees_din <= x"00a10801";
		wait for Clk_period;
		Addr <=  "00000111011101";
		Trees_din <= x"fff70801";
		wait for Clk_period;
		Addr <=  "00000111011110";
		Trees_din <= x"1400520c";
		wait for Clk_period;
		Addr <=  "00000111011111";
		Trees_din <= x"03fc9c08";
		wait for Clk_period;
		Addr <=  "00000111100000";
		Trees_din <= x"07005604";
		wait for Clk_period;
		Addr <=  "00000111100001";
		Trees_din <= x"00930801";
		wait for Clk_period;
		Addr <=  "00000111100010";
		Trees_din <= x"00210801";
		wait for Clk_period;
		Addr <=  "00000111100011";
		Trees_din <= x"ffb00801";
		wait for Clk_period;
		Addr <=  "00000111100100";
		Trees_din <= x"0b038f04";
		wait for Clk_period;
		Addr <=  "00000111100101";
		Trees_din <= x"ff7e0801";
		wait for Clk_period;
		Addr <=  "00000111100110";
		Trees_din <= x"fff50801";
		wait for Clk_period;
		Addr <=  "00000111100111";
		Trees_din <= x"050d5a1c";
		wait for Clk_period;
		Addr <=  "00000111101000";
		Trees_din <= x"020c5e18";
		wait for Clk_period;
		Addr <=  "00000111101001";
		Trees_din <= x"000e6e10";
		wait for Clk_period;
		Addr <=  "00000111101010";
		Trees_din <= x"0ef8d308";
		wait for Clk_period;
		Addr <=  "00000111101011";
		Trees_din <= x"0ef88004";
		wait for Clk_period;
		Addr <=  "00000111101100";
		Trees_din <= x"00120801";
		wait for Clk_period;
		Addr <=  "00000111101101";
		Trees_din <= x"ff830801";
		wait for Clk_period;
		Addr <=  "00000111101110";
		Trees_din <= x"02fa1e04";
		wait for Clk_period;
		Addr <=  "00000111101111";
		Trees_din <= x"ffa20801";
		wait for Clk_period;
		Addr <=  "00000111110000";
		Trees_din <= x"00660801";
		wait for Clk_period;
		Addr <=  "00000111110001";
		Trees_din <= x"1c004304";
		wait for Clk_period;
		Addr <=  "00000111110010";
		Trees_din <= x"ff870801";
		wait for Clk_period;
		Addr <=  "00000111110011";
		Trees_din <= x"00260801";
		wait for Clk_period;
		Addr <=  "00000111110100";
		Trees_din <= x"ff840801";
		wait for Clk_period;
		Addr <=  "00000111110101";
		Trees_din <= x"040ac910";
		wait for Clk_period;
		Addr <=  "00000111110110";
		Trees_din <= x"000b0b04";
		wait for Clk_period;
		Addr <=  "00000111110111";
		Trees_din <= x"00a40801";
		wait for Clk_period;
		Addr <=  "00000111111000";
		Trees_din <= x"06fc2004";
		wait for Clk_period;
		Addr <=  "00000111111001";
		Trees_din <= x"00920801";
		wait for Clk_period;
		Addr <=  "00000111111010";
		Trees_din <= x"03fcc704";
		wait for Clk_period;
		Addr <=  "00000111111011";
		Trees_din <= x"00440801";
		wait for Clk_period;
		Addr <=  "00000111111100";
		Trees_din <= x"ff8e0801";
		wait for Clk_period;
		Addr <=  "00000111111101";
		Trees_din <= x"0515e904";
		wait for Clk_period;
		Addr <=  "00000111111110";
		Trees_din <= x"ff930801";
		wait for Clk_period;
		Addr <=  "00000111111111";
		Trees_din <= x"00860801";
		wait for Clk_period;
		Addr <=  "00001000000000";
		Trees_din <= x"05085524";
		wait for Clk_period;
		Addr <=  "00001000000001";
		Trees_din <= x"0506f714";
		wait for Clk_period;
		Addr <=  "00001000000010";
		Trees_din <= x"20000e10";
		wait for Clk_period;
		Addr <=  "00001000000011";
		Trees_din <= x"0e017f04";
		wait for Clk_period;
		Addr <=  "00001000000100";
		Trees_din <= x"ff6608c5";
		wait for Clk_period;
		Addr <=  "00001000000101";
		Trees_din <= x"0b040208";
		wait for Clk_period;
		Addr <=  "00001000000110";
		Trees_din <= x"14000104";
		wait for Clk_period;
		Addr <=  "00001000000111";
		Trees_din <= x"002608c5";
		wait for Clk_period;
		Addr <=  "00001000001000";
		Trees_din <= x"ff7108c5";
		wait for Clk_period;
		Addr <=  "00001000001001";
		Trees_din <= x"008608c5";
		wait for Clk_period;
		Addr <=  "00001000001010";
		Trees_din <= x"fffe08c5";
		wait for Clk_period;
		Addr <=  "00001000001011";
		Trees_din <= x"14005208";
		wait for Clk_period;
		Addr <=  "00001000001100";
		Trees_din <= x"17004504";
		wait for Clk_period;
		Addr <=  "00001000001101";
		Trees_din <= x"ffd108c5";
		wait for Clk_period;
		Addr <=  "00001000001110";
		Trees_din <= x"006c08c5";
		wait for Clk_period;
		Addr <=  "00001000001111";
		Trees_din <= x"05081c04";
		wait for Clk_period;
		Addr <=  "00001000010000";
		Trees_din <= x"ff8608c5";
		wait for Clk_period;
		Addr <=  "00001000010001";
		Trees_din <= x"ffea08c5";
		wait for Clk_period;
		Addr <=  "00001000010010";
		Trees_din <= x"050d5a28";
		wait for Clk_period;
		Addr <=  "00001000010011";
		Trees_din <= x"03fcf110";
		wait for Clk_period;
		Addr <=  "00001000010100";
		Trees_din <= x"0208360c";
		wait for Clk_period;
		Addr <=  "00001000010101";
		Trees_din <= x"000b6404";
		wait for Clk_period;
		Addr <=  "00001000010110";
		Trees_din <= x"009808c5";
		wait for Clk_period;
		Addr <=  "00001000010111";
		Trees_din <= x"08005804";
		wait for Clk_period;
		Addr <=  "00001000011000";
		Trees_din <= x"ffd408c5";
		wait for Clk_period;
		Addr <=  "00001000011001";
		Trees_din <= x"008d08c5";
		wait for Clk_period;
		Addr <=  "00001000011010";
		Trees_din <= x"ffb508c5";
		wait for Clk_period;
		Addr <=  "00001000011011";
		Trees_din <= x"09f96b08";
		wait for Clk_period;
		Addr <=  "00001000011100";
		Trees_din <= x"1602dc04";
		wait for Clk_period;
		Addr <=  "00001000011101";
		Trees_din <= x"000208c5";
		wait for Clk_period;
		Addr <=  "00001000011110";
		Trees_din <= x"009a08c5";
		wait for Clk_period;
		Addr <=  "00001000011111";
		Trees_din <= x"000b0b08";
		wait for Clk_period;
		Addr <=  "00001000100000";
		Trees_din <= x"00ec0004";
		wait for Clk_period;
		Addr <=  "00001000100001";
		Trees_din <= x"ff8b08c5";
		wait for Clk_period;
		Addr <=  "00001000100010";
		Trees_din <= x"005c08c5";
		wait for Clk_period;
		Addr <=  "00001000100011";
		Trees_din <= x"1b034204";
		wait for Clk_period;
		Addr <=  "00001000100100";
		Trees_din <= x"ff7208c5";
		wait for Clk_period;
		Addr <=  "00001000100101";
		Trees_din <= x"ffe608c5";
		wait for Clk_period;
		Addr <=  "00001000100110";
		Trees_din <= x"040ac910";
		wait for Clk_period;
		Addr <=  "00001000100111";
		Trees_din <= x"000b0b04";
		wait for Clk_period;
		Addr <=  "00001000101000";
		Trees_din <= x"00a008c5";
		wait for Clk_period;
		Addr <=  "00001000101001";
		Trees_din <= x"1403ba08";
		wait for Clk_period;
		Addr <=  "00001000101010";
		Trees_din <= x"16000104";
		wait for Clk_period;
		Addr <=  "00001000101011";
		Trees_din <= x"ffe308c5";
		wait for Clk_period;
		Addr <=  "00001000101100";
		Trees_din <= x"008b08c5";
		wait for Clk_period;
		Addr <=  "00001000101101";
		Trees_din <= x"ffb408c5";
		wait for Clk_period;
		Addr <=  "00001000101110";
		Trees_din <= x"0515e904";
		wait for Clk_period;
		Addr <=  "00001000101111";
		Trees_din <= x"ff9b08c5";
		wait for Clk_period;
		Addr <=  "00001000110000";
		Trees_din <= x"007908c5";
		wait for Clk_period;
		Addr <=  "00001000110001";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00001000110010";
		Trees_din <= x"05081c20";
		wait for Clk_period;
		Addr <=  "00001000110011";
		Trees_din <= x"0506f714";
		wait for Clk_period;
		Addr <=  "00001000110100";
		Trees_din <= x"0e017f08";
		wait for Clk_period;
		Addr <=  "00001000110101";
		Trees_din <= x"20000e04";
		wait for Clk_period;
		Addr <=  "00001000110110";
		Trees_din <= x"ff670985";
		wait for Clk_period;
		Addr <=  "00001000110111";
		Trees_din <= x"000c0985";
		wait for Clk_period;
		Addr <=  "00001000111000";
		Trees_din <= x"0b040208";
		wait for Clk_period;
		Addr <=  "00001000111001";
		Trees_din <= x"18004e04";
		wait for Clk_period;
		Addr <=  "00001000111010";
		Trees_din <= x"ff740985";
		wait for Clk_period;
		Addr <=  "00001000111011";
		Trees_din <= x"00280985";
		wait for Clk_period;
		Addr <=  "00001000111100";
		Trees_din <= x"00780985";
		wait for Clk_period;
		Addr <=  "00001000111101";
		Trees_din <= x"0d03eb08";
		wait for Clk_period;
		Addr <=  "00001000111110";
		Trees_din <= x"16000004";
		wait for Clk_period;
		Addr <=  "00001000111111";
		Trees_din <= x"ffef0985";
		wait for Clk_period;
		Addr <=  "00001001000000";
		Trees_din <= x"ff8b0985";
		wait for Clk_period;
		Addr <=  "00001001000001";
		Trees_din <= x"00530985";
		wait for Clk_period;
		Addr <=  "00001001000010";
		Trees_din <= x"050d5a28";
		wait for Clk_period;
		Addr <=  "00001001000011";
		Trees_din <= x"00f45908";
		wait for Clk_period;
		Addr <=  "00001001000100";
		Trees_din <= x"03fd1f04";
		wait for Clk_period;
		Addr <=  "00001001000101";
		Trees_din <= x"fffb0985";
		wait for Clk_period;
		Addr <=  "00001001000110";
		Trees_din <= x"ff8b0985";
		wait for Clk_period;
		Addr <=  "00001001000111";
		Trees_din <= x"000b6410";
		wait for Clk_period;
		Addr <=  "00001001001000";
		Trees_din <= x"06fb1408";
		wait for Clk_period;
		Addr <=  "00001001001001";
		Trees_din <= x"12009e04";
		wait for Clk_period;
		Addr <=  "00001001001010";
		Trees_din <= x"00200985";
		wait for Clk_period;
		Addr <=  "00001001001011";
		Trees_din <= x"ffa80985";
		wait for Clk_period;
		Addr <=  "00001001001100";
		Trees_din <= x"11005304";
		wait for Clk_period;
		Addr <=  "00001001001101";
		Trees_din <= x"00270985";
		wait for Clk_period;
		Addr <=  "00001001001110";
		Trees_din <= x"00930985";
		wait for Clk_period;
		Addr <=  "00001001001111";
		Trees_din <= x"09fa5308";
		wait for Clk_period;
		Addr <=  "00001001010000";
		Trees_din <= x"08005304";
		wait for Clk_period;
		Addr <=  "00001001010001";
		Trees_din <= x"ffab0985";
		wait for Clk_period;
		Addr <=  "00001001010010";
		Trees_din <= x"00980985";
		wait for Clk_period;
		Addr <=  "00001001010011";
		Trees_din <= x"0904ad04";
		wait for Clk_period;
		Addr <=  "00001001010100";
		Trees_din <= x"ff880985";
		wait for Clk_period;
		Addr <=  "00001001010101";
		Trees_din <= x"00350985";
		wait for Clk_period;
		Addr <=  "00001001010110";
		Trees_din <= x"01184314";
		wait for Clk_period;
		Addr <=  "00001001010111";
		Trees_din <= x"000b0b08";
		wait for Clk_period;
		Addr <=  "00001001011000";
		Trees_din <= x"18005404";
		wait for Clk_period;
		Addr <=  "00001001011001";
		Trees_din <= x"009c0985";
		wait for Clk_period;
		Addr <=  "00001001011010";
		Trees_din <= x"00330985";
		wait for Clk_period;
		Addr <=  "00001001011011";
		Trees_din <= x"0d011b08";
		wait for Clk_period;
		Addr <=  "00001001011100";
		Trees_din <= x"0a001404";
		wait for Clk_period;
		Addr <=  "00001001011101";
		Trees_din <= x"005e0985";
		wait for Clk_period;
		Addr <=  "00001001011110";
		Trees_din <= x"ffa50985";
		wait for Clk_period;
		Addr <=  "00001001011111";
		Trees_din <= x"007f0985";
		wait for Clk_period;
		Addr <=  "00001001100000";
		Trees_din <= x"fff50985";
		wait for Clk_period;
		Addr <=  "00001001100001";
		Trees_din <= x"05081c20";
		wait for Clk_period;
		Addr <=  "00001001100010";
		Trees_din <= x"18004e14";
		wait for Clk_period;
		Addr <=  "00001001100011";
		Trees_din <= x"0b04020c";
		wait for Clk_period;
		Addr <=  "00001001100100";
		Trees_din <= x"04fd7604";
		wait for Clk_period;
		Addr <=  "00001001100101";
		Trees_din <= x"fff30a49";
		wait for Clk_period;
		Addr <=  "00001001100110";
		Trees_din <= x"03fa1004";
		wait for Clk_period;
		Addr <=  "00001001100111";
		Trees_din <= x"ffc90a49";
		wait for Clk_period;
		Addr <=  "00001001101000";
		Trees_din <= x"ff680a49";
		wait for Clk_period;
		Addr <=  "00001001101001";
		Trees_din <= x"0e017f04";
		wait for Clk_period;
		Addr <=  "00001001101010";
		Trees_din <= x"ff800a49";
		wait for Clk_period;
		Addr <=  "00001001101011";
		Trees_din <= x"00670a49";
		wait for Clk_period;
		Addr <=  "00001001101100";
		Trees_din <= x"03fd0f08";
		wait for Clk_period;
		Addr <=  "00001001101101";
		Trees_din <= x"0d035d04";
		wait for Clk_period;
		Addr <=  "00001001101110";
		Trees_din <= x"00070a49";
		wait for Clk_period;
		Addr <=  "00001001101111";
		Trees_din <= x"00820a49";
		wait for Clk_period;
		Addr <=  "00001001110000";
		Trees_din <= x"ff880a49";
		wait for Clk_period;
		Addr <=  "00001001110001";
		Trees_din <= x"050d5a2c";
		wait for Clk_period;
		Addr <=  "00001001110010";
		Trees_din <= x"03fcf114";
		wait for Clk_period;
		Addr <=  "00001001110011";
		Trees_din <= x"08004e08";
		wait for Clk_period;
		Addr <=  "00001001110100";
		Trees_din <= x"050a6c04";
		wait for Clk_period;
		Addr <=  "00001001110101";
		Trees_din <= x"ff9e0a49";
		wait for Clk_period;
		Addr <=  "00001001110110";
		Trees_din <= x"00150a49";
		wait for Clk_period;
		Addr <=  "00001001110111";
		Trees_din <= x"0ef8ee04";
		wait for Clk_period;
		Addr <=  "00001001111000";
		Trees_din <= x"ffca0a49";
		wait for Clk_period;
		Addr <=  "00001001111001";
		Trees_din <= x"0c018d04";
		wait for Clk_period;
		Addr <=  "00001001111010";
		Trees_din <= x"00820a49";
		wait for Clk_period;
		Addr <=  "00001001111011";
		Trees_din <= x"001a0a49";
		wait for Clk_period;
		Addr <=  "00001001111100";
		Trees_din <= x"04fe0d0c";
		wait for Clk_period;
		Addr <=  "00001001111101";
		Trees_din <= x"0efedf04";
		wait for Clk_period;
		Addr <=  "00001001111110";
		Trees_din <= x"ffcf0a49";
		wait for Clk_period;
		Addr <=  "00001001111111";
		Trees_din <= x"08005604";
		wait for Clk_period;
		Addr <=  "00001010000000";
		Trees_din <= x"00090a49";
		wait for Clk_period;
		Addr <=  "00001010000001";
		Trees_din <= x"008b0a49";
		wait for Clk_period;
		Addr <=  "00001010000010";
		Trees_din <= x"0c02c208";
		wait for Clk_period;
		Addr <=  "00001010000011";
		Trees_din <= x"0c008504";
		wait for Clk_period;
		Addr <=  "00001010000100";
		Trees_din <= x"fff20a49";
		wait for Clk_period;
		Addr <=  "00001010000101";
		Trees_din <= x"ff850a49";
		wait for Clk_period;
		Addr <=  "00001010000110";
		Trees_din <= x"00260a49";
		wait for Clk_period;
		Addr <=  "00001010000111";
		Trees_din <= x"040ac910";
		wait for Clk_period;
		Addr <=  "00001010001000";
		Trees_din <= x"000b0b04";
		wait for Clk_period;
		Addr <=  "00001010001001";
		Trees_din <= x"00990a49";
		wait for Clk_period;
		Addr <=  "00001010001010";
		Trees_din <= x"0b02cb08";
		wait for Clk_period;
		Addr <=  "00001010001011";
		Trees_din <= x"03fcc704";
		wait for Clk_period;
		Addr <=  "00001010001100";
		Trees_din <= x"00840a49";
		wait for Clk_period;
		Addr <=  "00001010001101";
		Trees_din <= x"fffe0a49";
		wait for Clk_period;
		Addr <=  "00001010001110";
		Trees_din <= x"ffc70a49";
		wait for Clk_period;
		Addr <=  "00001010001111";
		Trees_din <= x"051b3b04";
		wait for Clk_period;
		Addr <=  "00001010010000";
		Trees_din <= x"ffb70a49";
		wait for Clk_period;
		Addr <=  "00001010010001";
		Trees_din <= x"00770a49";
		wait for Clk_period;
		Addr <=  "00001010010010";
		Trees_din <= x"05072418";
		wait for Clk_period;
		Addr <=  "00001010010011";
		Trees_din <= x"0e017f0c";
		wait for Clk_period;
		Addr <=  "00001010010100";
		Trees_din <= x"03fac208";
		wait for Clk_period;
		Addr <=  "00001010010101";
		Trees_din <= x"05052c04";
		wait for Clk_period;
		Addr <=  "00001010010110";
		Trees_din <= x"ffa20b05";
		wait for Clk_period;
		Addr <=  "00001010010111";
		Trees_din <= x"00430b05";
		wait for Clk_period;
		Addr <=  "00001010011000";
		Trees_din <= x"ff690b05";
		wait for Clk_period;
		Addr <=  "00001010011001";
		Trees_din <= x"0e018704";
		wait for Clk_period;
		Addr <=  "00001010011010";
		Trees_din <= x"00690b05";
		wait for Clk_period;
		Addr <=  "00001010011011";
		Trees_din <= x"08005904";
		wait for Clk_period;
		Addr <=  "00001010011100";
		Trees_din <= x"ff7e0b05";
		wait for Clk_period;
		Addr <=  "00001010011101";
		Trees_din <= x"00140b05";
		wait for Clk_period;
		Addr <=  "00001010011110";
		Trees_din <= x"050d5a30";
		wait for Clk_period;
		Addr <=  "00001010011111";
		Trees_din <= x"03fcf11c";
		wait for Clk_period;
		Addr <=  "00001010100000";
		Trees_din <= x"0a013b10";
		wait for Clk_period;
		Addr <=  "00001010100001";
		Trees_din <= x"0904a908";
		wait for Clk_period;
		Addr <=  "00001010100010";
		Trees_din <= x"000a8004";
		wait for Clk_period;
		Addr <=  "00001010100011";
		Trees_din <= x"00110b05";
		wait for Clk_period;
		Addr <=  "00001010100100";
		Trees_din <= x"ff840b05";
		wait for Clk_period;
		Addr <=  "00001010100101";
		Trees_din <= x"0c008304";
		wait for Clk_period;
		Addr <=  "00001010100110";
		Trees_din <= x"006b0b05";
		wait for Clk_period;
		Addr <=  "00001010100111";
		Trees_din <= x"fffe0b05";
		wait for Clk_period;
		Addr <=  "00001010101000";
		Trees_din <= x"12009404";
		wait for Clk_period;
		Addr <=  "00001010101001";
		Trees_din <= x"009e0b05";
		wait for Clk_period;
		Addr <=  "00001010101010";
		Trees_din <= x"000b6404";
		wait for Clk_period;
		Addr <=  "00001010101011";
		Trees_din <= x"00410b05";
		wait for Clk_period;
		Addr <=  "00001010101100";
		Trees_din <= x"ffca0b05";
		wait for Clk_period;
		Addr <=  "00001010101101";
		Trees_din <= x"09f96b04";
		wait for Clk_period;
		Addr <=  "00001010101110";
		Trees_din <= x"00460b05";
		wait for Clk_period;
		Addr <=  "00001010101111";
		Trees_din <= x"000b0b08";
		wait for Clk_period;
		Addr <=  "00001010110000";
		Trees_din <= x"00ec0004";
		wait for Clk_period;
		Addr <=  "00001010110001";
		Trees_din <= x"ff980b05";
		wait for Clk_period;
		Addr <=  "00001010110010";
		Trees_din <= x"00440b05";
		wait for Clk_period;
		Addr <=  "00001010110011";
		Trees_din <= x"16000004";
		wait for Clk_period;
		Addr <=  "00001010110100";
		Trees_din <= x"ffdc0b05";
		wait for Clk_period;
		Addr <=  "00001010110101";
		Trees_din <= x"ff7f0b05";
		wait for Clk_period;
		Addr <=  "00001010110110";
		Trees_din <= x"040ac910";
		wait for Clk_period;
		Addr <=  "00001010110111";
		Trees_din <= x"000b0b04";
		wait for Clk_period;
		Addr <=  "00001010111000";
		Trees_din <= x"00960b05";
		wait for Clk_period;
		Addr <=  "00001010111001";
		Trees_din <= x"06fc2004";
		wait for Clk_period;
		Addr <=  "00001010111010";
		Trees_din <= x"006e0b05";
		wait for Clk_period;
		Addr <=  "00001010111011";
		Trees_din <= x"01f96404";
		wait for Clk_period;
		Addr <=  "00001010111100";
		Trees_din <= x"ffa80b05";
		wait for Clk_period;
		Addr <=  "00001010111101";
		Trees_din <= x"00320b05";
		wait for Clk_period;
		Addr <=  "00001010111110";
		Trees_din <= x"0515e904";
		wait for Clk_period;
		Addr <=  "00001010111111";
		Trees_din <= x"ffab0b05";
		wait for Clk_period;
		Addr <=  "00001011000000";
		Trees_din <= x"00600b05";
		wait for Clk_period;
		Addr <=  "00001011000001";
		Trees_din <= x"05072418";
		wait for Clk_period;
		Addr <=  "00001011000010";
		Trees_din <= x"0e017f0c";
		wait for Clk_period;
		Addr <=  "00001011000011";
		Trees_din <= x"03fac208";
		wait for Clk_period;
		Addr <=  "00001011000100";
		Trees_din <= x"05052c04";
		wait for Clk_period;
		Addr <=  "00001011000101";
		Trees_din <= x"ffa90b99";
		wait for Clk_period;
		Addr <=  "00001011000110";
		Trees_din <= x"003a0b99";
		wait for Clk_period;
		Addr <=  "00001011000111";
		Trees_din <= x"ff6a0b99";
		wait for Clk_period;
		Addr <=  "00001011001000";
		Trees_din <= x"0b040208";
		wait for Clk_period;
		Addr <=  "00001011001001";
		Trees_din <= x"19007b04";
		wait for Clk_period;
		Addr <=  "00001011001010";
		Trees_din <= x"00100b99";
		wait for Clk_period;
		Addr <=  "00001011001011";
		Trees_din <= x"ff840b99";
		wait for Clk_period;
		Addr <=  "00001011001100";
		Trees_din <= x"00640b99";
		wait for Clk_period;
		Addr <=  "00001011001101";
		Trees_din <= x"0510932c";
		wait for Clk_period;
		Addr <=  "00001011001110";
		Trees_din <= x"03fcf114";
		wait for Clk_period;
		Addr <=  "00001011001111";
		Trees_din <= x"1403ee0c";
		wait for Clk_period;
		Addr <=  "00001011010000";
		Trees_din <= x"020b1e08";
		wait for Clk_period;
		Addr <=  "00001011010001";
		Trees_din <= x"000b6404";
		wait for Clk_period;
		Addr <=  "00001011010010";
		Trees_din <= x"008b0b99";
		wait for Clk_period;
		Addr <=  "00001011010011";
		Trees_din <= x"003a0b99";
		wait for Clk_period;
		Addr <=  "00001011010100";
		Trees_din <= x"ffdb0b99";
		wait for Clk_period;
		Addr <=  "00001011010101";
		Trees_din <= x"07005804";
		wait for Clk_period;
		Addr <=  "00001011010110";
		Trees_din <= x"000d0b99";
		wait for Clk_period;
		Addr <=  "00001011010111";
		Trees_din <= x"ffbd0b99";
		wait for Clk_period;
		Addr <=  "00001011011000";
		Trees_din <= x"04feaa0c";
		wait for Clk_period;
		Addr <=  "00001011011001";
		Trees_din <= x"000b0b04";
		wait for Clk_period;
		Addr <=  "00001011011010";
		Trees_din <= x"00670b99";
		wait for Clk_period;
		Addr <=  "00001011011011";
		Trees_din <= x"09f96b04";
		wait for Clk_period;
		Addr <=  "00001011011100";
		Trees_din <= x"005b0b99";
		wait for Clk_period;
		Addr <=  "00001011011101";
		Trees_din <= x"ffb40b99";
		wait for Clk_period;
		Addr <=  "00001011011110";
		Trees_din <= x"0c029608";
		wait for Clk_period;
		Addr <=  "00001011011111";
		Trees_din <= x"0c004504";
		wait for Clk_period;
		Addr <=  "00001011100000";
		Trees_din <= x"ffeb0b99";
		wait for Clk_period;
		Addr <=  "00001011100001";
		Trees_din <= x"ff920b99";
		wait for Clk_period;
		Addr <=  "00001011100010";
		Trees_din <= x"00200b99";
		wait for Clk_period;
		Addr <=  "00001011100011";
		Trees_din <= x"03092d04";
		wait for Clk_period;
		Addr <=  "00001011100100";
		Trees_din <= x"00980b99";
		wait for Clk_period;
		Addr <=  "00001011100101";
		Trees_din <= x"00210b99";
		wait for Clk_period;
		Addr <=  "00001011100110";
		Trees_din <= x"05085518";
		wait for Clk_period;
		Addr <=  "00001011100111";
		Trees_din <= x"05039508";
		wait for Clk_period;
		Addr <=  "00001011101000";
		Trees_din <= x"15f8e904";
		wait for Clk_period;
		Addr <=  "00001011101001";
		Trees_din <= x"001c0c15";
		wait for Clk_period;
		Addr <=  "00001011101010";
		Trees_din <= x"ff6b0c15";
		wait for Clk_period;
		Addr <=  "00001011101011";
		Trees_din <= x"18004e0c";
		wait for Clk_period;
		Addr <=  "00001011101100";
		Trees_din <= x"0a02fb04";
		wait for Clk_period;
		Addr <=  "00001011101101";
		Trees_din <= x"ff850c15";
		wait for Clk_period;
		Addr <=  "00001011101110";
		Trees_din <= x"01fd5304";
		wait for Clk_period;
		Addr <=  "00001011101111";
		Trees_din <= x"ffa80c15";
		wait for Clk_period;
		Addr <=  "00001011110000";
		Trees_din <= x"00380c15";
		wait for Clk_period;
		Addr <=  "00001011110001";
		Trees_din <= x"00450c15";
		wait for Clk_period;
		Addr <=  "00001011110010";
		Trees_din <= x"05109320";
		wait for Clk_period;
		Addr <=  "00001011110011";
		Trees_din <= x"020e161c";
		wait for Clk_period;
		Addr <=  "00001011110100";
		Trees_din <= x"08005210";
		wait for Clk_period;
		Addr <=  "00001011110101";
		Trees_din <= x"01fa2a08";
		wait for Clk_period;
		Addr <=  "00001011110110";
		Trees_din <= x"19009404";
		wait for Clk_period;
		Addr <=  "00001011110111";
		Trees_din <= x"fff50c15";
		wait for Clk_period;
		Addr <=  "00001011111000";
		Trees_din <= x"ffa10c15";
		wait for Clk_period;
		Addr <=  "00001011111001";
		Trees_din <= x"0509dd04";
		wait for Clk_period;
		Addr <=  "00001011111010";
		Trees_din <= x"ffd20c15";
		wait for Clk_period;
		Addr <=  "00001011111011";
		Trees_din <= x"00540c15";
		wait for Clk_period;
		Addr <=  "00001011111100";
		Trees_din <= x"02fa3b04";
		wait for Clk_period;
		Addr <=  "00001011111101";
		Trees_din <= x"ffd30c15";
		wait for Clk_period;
		Addr <=  "00001011111110";
		Trees_din <= x"11039a04";
		wait for Clk_period;
		Addr <=  "00001011111111";
		Trees_din <= x"006f0c15";
		wait for Clk_period;
		Addr <=  "00001100000000";
		Trees_din <= x"00070c15";
		wait for Clk_period;
		Addr <=  "00001100000001";
		Trees_din <= x"ff9c0c15";
		wait for Clk_period;
		Addr <=  "00001100000010";
		Trees_din <= x"03092d04";
		wait for Clk_period;
		Addr <=  "00001100000011";
		Trees_din <= x"00960c15";
		wait for Clk_period;
		Addr <=  "00001100000100";
		Trees_din <= x"00210c15";
		wait for Clk_period;
		Addr <=  "00001100000101";
		Trees_din <= x"05072414";
		wait for Clk_period;
		Addr <=  "00001100000110";
		Trees_din <= x"0e017f08";
		wait for Clk_period;
		Addr <=  "00001100000111";
		Trees_din <= x"03fac204";
		wait for Clk_period;
		Addr <=  "00001100001000";
		Trees_din <= x"ffef0c99";
		wait for Clk_period;
		Addr <=  "00001100001001";
		Trees_din <= x"ff6d0c99";
		wait for Clk_period;
		Addr <=  "00001100001010";
		Trees_din <= x"0e018704";
		wait for Clk_period;
		Addr <=  "00001100001011";
		Trees_din <= x"00690c99";
		wait for Clk_period;
		Addr <=  "00001100001100";
		Trees_din <= x"0c005104";
		wait for Clk_period;
		Addr <=  "00001100001101";
		Trees_din <= x"00020c99";
		wait for Clk_period;
		Addr <=  "00001100001110";
		Trees_din <= x"ff930c99";
		wait for Clk_period;
		Addr <=  "00001100001111";
		Trees_din <= x"050d5a18";
		wait for Clk_period;
		Addr <=  "00001100010000";
		Trees_din <= x"0ef8f704";
		wait for Clk_period;
		Addr <=  "00001100010001";
		Trees_din <= x"ffad0c99";
		wait for Clk_period;
		Addr <=  "00001100010010";
		Trees_din <= x"01027c10";
		wait for Clk_period;
		Addr <=  "00001100010011";
		Trees_din <= x"01fa7a08";
		wait for Clk_period;
		Addr <=  "00001100010100";
		Trees_din <= x"0c00ba04";
		wait for Clk_period;
		Addr <=  "00001100010101";
		Trees_din <= x"00370c99";
		wait for Clk_period;
		Addr <=  "00001100010110";
		Trees_din <= x"ffaf0c99";
		wait for Clk_period;
		Addr <=  "00001100010111";
		Trees_din <= x"0b03c004";
		wait for Clk_period;
		Addr <=  "00001100011000";
		Trees_din <= x"005f0c99";
		wait for Clk_period;
		Addr <=  "00001100011001";
		Trees_din <= x"ffe20c99";
		wait for Clk_period;
		Addr <=  "00001100011010";
		Trees_din <= x"ffb20c99";
		wait for Clk_period;
		Addr <=  "00001100011011";
		Trees_din <= x"040ac910";
		wait for Clk_period;
		Addr <=  "00001100011100";
		Trees_din <= x"000b0b04";
		wait for Clk_period;
		Addr <=  "00001100011101";
		Trees_din <= x"008f0c99";
		wait for Clk_period;
		Addr <=  "00001100011110";
		Trees_din <= x"050f3508";
		wait for Clk_period;
		Addr <=  "00001100011111";
		Trees_din <= x"1300fe04";
		wait for Clk_period;
		Addr <=  "00001100100000";
		Trees_din <= x"00620c99";
		wait for Clk_period;
		Addr <=  "00001100100001";
		Trees_din <= x"00190c99";
		wait for Clk_period;
		Addr <=  "00001100100010";
		Trees_din <= x"ffdf0c99";
		wait for Clk_period;
		Addr <=  "00001100100011";
		Trees_din <= x"14015b04";
		wait for Clk_period;
		Addr <=  "00001100100100";
		Trees_din <= x"00510c99";
		wait for Clk_period;
		Addr <=  "00001100100101";
		Trees_din <= x"ffc10c99";
		wait for Clk_period;
		Addr <=  "00001100100110";
		Trees_din <= x"05081c18";
		wait for Clk_period;
		Addr <=  "00001100100111";
		Trees_din <= x"0e017f0c";
		wait for Clk_period;
		Addr <=  "00001100101000";
		Trees_din <= x"03fbcb08";
		wait for Clk_period;
		Addr <=  "00001100101001";
		Trees_din <= x"05054b04";
		wait for Clk_period;
		Addr <=  "00001100101010";
		Trees_din <= x"ffa10d1d";
		wait for Clk_period;
		Addr <=  "00001100101011";
		Trees_din <= x"00330d1d";
		wait for Clk_period;
		Addr <=  "00001100101100";
		Trees_din <= x"ff700d1d";
		wait for Clk_period;
		Addr <=  "00001100101101";
		Trees_din <= x"0b040208";
		wait for Clk_period;
		Addr <=  "00001100101110";
		Trees_din <= x"03fd0f04";
		wait for Clk_period;
		Addr <=  "00001100101111";
		Trees_din <= x"00000d1d";
		wait for Clk_period;
		Addr <=  "00001100110000";
		Trees_din <= x"ff9a0d1d";
		wait for Clk_period;
		Addr <=  "00001100110001";
		Trees_din <= x"005d0d1d";
		wait for Clk_period;
		Addr <=  "00001100110010";
		Trees_din <= x"05109324";
		wait for Clk_period;
		Addr <=  "00001100110011";
		Trees_din <= x"00f1de08";
		wait for Clk_period;
		Addr <=  "00001100110100";
		Trees_din <= x"0403e804";
		wait for Clk_period;
		Addr <=  "00001100110101";
		Trees_din <= x"fff20d1d";
		wait for Clk_period;
		Addr <=  "00001100110110";
		Trees_din <= x"ffa50d1d";
		wait for Clk_period;
		Addr <=  "00001100110111";
		Trees_din <= x"000b0b0c";
		wait for Clk_period;
		Addr <=  "00001100111000";
		Trees_din <= x"02088f08";
		wait for Clk_period;
		Addr <=  "00001100111001";
		Trees_din <= x"1d00f304";
		wait for Clk_period;
		Addr <=  "00001100111010";
		Trees_din <= x"00830d1d";
		wait for Clk_period;
		Addr <=  "00001100111011";
		Trees_din <= x"00120d1d";
		wait for Clk_period;
		Addr <=  "00001100111100";
		Trees_din <= x"fff80d1d";
		wait for Clk_period;
		Addr <=  "00001100111101";
		Trees_din <= x"0a013b08";
		wait for Clk_period;
		Addr <=  "00001100111110";
		Trees_din <= x"13fafb04";
		wait for Clk_period;
		Addr <=  "00001100111111";
		Trees_din <= x"00350d1d";
		wait for Clk_period;
		Addr <=  "00001101000000";
		Trees_din <= x"ffb10d1d";
		wait for Clk_period;
		Addr <=  "00001101000001";
		Trees_din <= x"01fa0c04";
		wait for Clk_period;
		Addr <=  "00001101000010";
		Trees_din <= x"ffda0d1d";
		wait for Clk_period;
		Addr <=  "00001101000011";
		Trees_din <= x"005e0d1d";
		wait for Clk_period;
		Addr <=  "00001101000100";
		Trees_din <= x"03092d04";
		wait for Clk_period;
		Addr <=  "00001101000101";
		Trees_din <= x"00900d1d";
		wait for Clk_period;
		Addr <=  "00001101000110";
		Trees_din <= x"001c0d1d";
		wait for Clk_period;
		Addr <=  "00001101000111";
		Trees_din <= x"05085518";
		wait for Clk_period;
		Addr <=  "00001101001000";
		Trees_din <= x"0e017f0c";
		wait for Clk_period;
		Addr <=  "00001101001001";
		Trees_din <= x"05054b04";
		wait for Clk_period;
		Addr <=  "00001101001010";
		Trees_din <= x"ff710d99";
		wait for Clk_period;
		Addr <=  "00001101001011";
		Trees_din <= x"03fbcb04";
		wait for Clk_period;
		Addr <=  "00001101001100";
		Trees_din <= x"00290d99";
		wait for Clk_period;
		Addr <=  "00001101001101";
		Trees_din <= x"ffac0d99";
		wait for Clk_period;
		Addr <=  "00001101001110";
		Trees_din <= x"000b0b08";
		wait for Clk_period;
		Addr <=  "00001101001111";
		Trees_din <= x"02ffab04";
		wait for Clk_period;
		Addr <=  "00001101010000";
		Trees_din <= x"007c0d99";
		wait for Clk_period;
		Addr <=  "00001101010001";
		Trees_din <= x"ffe90d99";
		wait for Clk_period;
		Addr <=  "00001101010010";
		Trees_din <= x"ffa10d99";
		wait for Clk_period;
		Addr <=  "00001101010011";
		Trees_din <= x"05109320";
		wait for Clk_period;
		Addr <=  "00001101010100";
		Trees_din <= x"020e161c";
		wait for Clk_period;
		Addr <=  "00001101010101";
		Trees_din <= x"0800520c";
		wait for Clk_period;
		Addr <=  "00001101010110";
		Trees_din <= x"0c002104";
		wait for Clk_period;
		Addr <=  "00001101010111";
		Trees_din <= x"00530d99";
		wait for Clk_period;
		Addr <=  "00001101011000";
		Trees_din <= x"00087604";
		wait for Clk_period;
		Addr <=  "00001101011001";
		Trees_din <= x"001f0d99";
		wait for Clk_period;
		Addr <=  "00001101011010";
		Trees_din <= x"ffae0d99";
		wait for Clk_period;
		Addr <=  "00001101011011";
		Trees_din <= x"04fecb08";
		wait for Clk_period;
		Addr <=  "00001101011100";
		Trees_din <= x"10021e04";
		wait for Clk_period;
		Addr <=  "00001101011101";
		Trees_din <= x"006e0d99";
		wait for Clk_period;
		Addr <=  "00001101011110";
		Trees_din <= x"00150d99";
		wait for Clk_period;
		Addr <=  "00001101011111";
		Trees_din <= x"11027a04";
		wait for Clk_period;
		Addr <=  "00001101100000";
		Trees_din <= x"00300d99";
		wait for Clk_period;
		Addr <=  "00001101100001";
		Trees_din <= x"ffbb0d99";
		wait for Clk_period;
		Addr <=  "00001101100010";
		Trees_din <= x"ffaa0d99";
		wait for Clk_period;
		Addr <=  "00001101100011";
		Trees_din <= x"03092d04";
		wait for Clk_period;
		Addr <=  "00001101100100";
		Trees_din <= x"008d0d99";
		wait for Clk_period;
		Addr <=  "00001101100101";
		Trees_din <= x"001b0d99";
		wait for Clk_period;
		Addr <=  "00001101100110";
		Trees_din <= x"05085518";
		wait for Clk_period;
		Addr <=  "00001101100111";
		Trees_din <= x"0e017f0c";
		wait for Clk_period;
		Addr <=  "00001101101000";
		Trees_din <= x"05054b04";
		wait for Clk_period;
		Addr <=  "00001101101001";
		Trees_din <= x"ff740e25";
		wait for Clk_period;
		Addr <=  "00001101101010";
		Trees_din <= x"12008404";
		wait for Clk_period;
		Addr <=  "00001101101011";
		Trees_din <= x"002d0e25";
		wait for Clk_period;
		Addr <=  "00001101101100";
		Trees_din <= x"ffb80e25";
		wait for Clk_period;
		Addr <=  "00001101101101";
		Trees_din <= x"000b0b08";
		wait for Clk_period;
		Addr <=  "00001101101110";
		Trees_din <= x"02ffab04";
		wait for Clk_period;
		Addr <=  "00001101101111";
		Trees_din <= x"006b0e25";
		wait for Clk_period;
		Addr <=  "00001101110000";
		Trees_din <= x"ffed0e25";
		wait for Clk_period;
		Addr <=  "00001101110001";
		Trees_din <= x"ffa90e25";
		wait for Clk_period;
		Addr <=  "00001101110010";
		Trees_din <= x"05109328";
		wait for Clk_period;
		Addr <=  "00001101110011";
		Trees_din <= x"03fcf114";
		wait for Clk_period;
		Addr <=  "00001101110100";
		Trees_din <= x"08005108";
		wait for Clk_period;
		Addr <=  "00001101110101";
		Trees_din <= x"07005604";
		wait for Clk_period;
		Addr <=  "00001101110110";
		Trees_din <= x"002b0e25";
		wait for Clk_period;
		Addr <=  "00001101110111";
		Trees_din <= x"ffbd0e25";
		wait for Clk_period;
		Addr <=  "00001101111000";
		Trees_din <= x"06fcf608";
		wait for Clk_period;
		Addr <=  "00001101111001";
		Trees_din <= x"000c1004";
		wait for Clk_period;
		Addr <=  "00001101111010";
		Trees_din <= x"004d0e25";
		wait for Clk_period;
		Addr <=  "00001101111011";
		Trees_din <= x"ffee0e25";
		wait for Clk_period;
		Addr <=  "00001101111100";
		Trees_din <= x"00750e25";
		wait for Clk_period;
		Addr <=  "00001101111101";
		Trees_din <= x"06fc2008";
		wait for Clk_period;
		Addr <=  "00001101111110";
		Trees_din <= x"1c003804";
		wait for Clk_period;
		Addr <=  "00001101111111";
		Trees_din <= x"ffee0e25";
		wait for Clk_period;
		Addr <=  "00001110000000";
		Trees_din <= x"004e0e25";
		wait for Clk_period;
		Addr <=  "00001110000001";
		Trees_din <= x"000b0b08";
		wait for Clk_period;
		Addr <=  "00001110000010";
		Trees_din <= x"00e9ab04";
		wait for Clk_period;
		Addr <=  "00001110000011";
		Trees_din <= x"ffbb0e25";
		wait for Clk_period;
		Addr <=  "00001110000100";
		Trees_din <= x"00490e25";
		wait for Clk_period;
		Addr <=  "00001110000101";
		Trees_din <= x"ffa70e25";
		wait for Clk_period;
		Addr <=  "00001110000110";
		Trees_din <= x"03092d04";
		wait for Clk_period;
		Addr <=  "00001110000111";
		Trees_din <= x"00890e25";
		wait for Clk_period;
		Addr <=  "00001110001000";
		Trees_din <= x"001a0e25";
		wait for Clk_period;
		Addr <=  "00001110001001";
		Trees_din <= x"05085518";
		wait for Clk_period;
		Addr <=  "00001110001010";
		Trees_din <= x"0e017f0c";
		wait for Clk_period;
		Addr <=  "00001110001011";
		Trees_din <= x"05054b04";
		wait for Clk_period;
		Addr <=  "00001110001100";
		Trees_din <= x"ff780eb1";
		wait for Clk_period;
		Addr <=  "00001110001101";
		Trees_din <= x"03fbcb04";
		wait for Clk_period;
		Addr <=  "00001110001110";
		Trees_din <= x"00220eb1";
		wait for Clk_period;
		Addr <=  "00001110001111";
		Trees_din <= x"ffb70eb1";
		wait for Clk_period;
		Addr <=  "00001110010000";
		Trees_din <= x"06ff1b04";
		wait for Clk_period;
		Addr <=  "00001110010001";
		Trees_din <= x"ffb10eb1";
		wait for Clk_period;
		Addr <=  "00001110010010";
		Trees_din <= x"03fdbf04";
		wait for Clk_period;
		Addr <=  "00001110010011";
		Trees_din <= x"00610eb1";
		wait for Clk_period;
		Addr <=  "00001110010100";
		Trees_din <= x"ffeb0eb1";
		wait for Clk_period;
		Addr <=  "00001110010101";
		Trees_din <= x"050d5a20";
		wait for Clk_period;
		Addr <=  "00001110010110";
		Trees_din <= x"0800540c";
		wait for Clk_period;
		Addr <=  "00001110010111";
		Trees_din <= x"09050808";
		wait for Clk_period;
		Addr <=  "00001110011000";
		Trees_din <= x"0f027304";
		wait for Clk_period;
		Addr <=  "00001110011001";
		Trees_din <= x"ffa10eb1";
		wait for Clk_period;
		Addr <=  "00001110011010";
		Trees_din <= x"00020eb1";
		wait for Clk_period;
		Addr <=  "00001110011011";
		Trees_din <= x"00320eb1";
		wait for Clk_period;
		Addr <=  "00001110011100";
		Trees_din <= x"02fde808";
		wait for Clk_period;
		Addr <=  "00001110011101";
		Trees_din <= x"1b019004";
		wait for Clk_period;
		Addr <=  "00001110011110";
		Trees_din <= x"00160eb1";
		wait for Clk_period;
		Addr <=  "00001110011111";
		Trees_din <= x"ffb40eb1";
		wait for Clk_period;
		Addr <=  "00001110100000";
		Trees_din <= x"04fda904";
		wait for Clk_period;
		Addr <=  "00001110100001";
		Trees_din <= x"ffe50eb1";
		wait for Clk_period;
		Addr <=  "00001110100010";
		Trees_din <= x"02002b04";
		wait for Clk_period;
		Addr <=  "00001110100011";
		Trees_din <= x"00740eb1";
		wait for Clk_period;
		Addr <=  "00001110100100";
		Trees_din <= x"00240eb1";
		wait for Clk_period;
		Addr <=  "00001110100101";
		Trees_din <= x"0308690c";
		wait for Clk_period;
		Addr <=  "00001110100110";
		Trees_din <= x"000b0b04";
		wait for Clk_period;
		Addr <=  "00001110100111";
		Trees_din <= x"007d0eb1";
		wait for Clk_period;
		Addr <=  "00001110101000";
		Trees_din <= x"06fc2004";
		wait for Clk_period;
		Addr <=  "00001110101001";
		Trees_din <= x"004a0eb1";
		wait for Clk_period;
		Addr <=  "00001110101010";
		Trees_din <= x"ffee0eb1";
		wait for Clk_period;
		Addr <=  "00001110101011";
		Trees_din <= x"00100eb1";
		wait for Clk_period;
		Addr <=  "00001110101100";
		Trees_din <= x"0506f70c";
		wait for Clk_period;
		Addr <=  "00001110101101";
		Trees_din <= x"0e017f04";
		wait for Clk_period;
		Addr <=  "00001110101110";
		Trees_din <= x"ff820f25";
		wait for Clk_period;
		Addr <=  "00001110101111";
		Trees_din <= x"0e018704";
		wait for Clk_period;
		Addr <=  "00001110110000";
		Trees_din <= x"00480f25";
		wait for Clk_period;
		Addr <=  "00001110110001";
		Trees_din <= x"ffcd0f25";
		wait for Clk_period;
		Addr <=  "00001110110010";
		Trees_din <= x"0510932c";
		wait for Clk_period;
		Addr <=  "00001110110011";
		Trees_din <= x"03fcf118";
		wait for Clk_period;
		Addr <=  "00001110110100";
		Trees_din <= x"0a013b0c";
		wait for Clk_period;
		Addr <=  "00001110110101";
		Trees_din <= x"050c4e08";
		wait for Clk_period;
		Addr <=  "00001110110110";
		Trees_din <= x"0c008704";
		wait for Clk_period;
		Addr <=  "00001110110111";
		Trees_din <= x"fffa0f25";
		wait for Clk_period;
		Addr <=  "00001110111000";
		Trees_din <= x"ffb40f25";
		wait for Clk_period;
		Addr <=  "00001110111001";
		Trees_din <= x"00460f25";
		wait for Clk_period;
		Addr <=  "00001110111010";
		Trees_din <= x"12009404";
		wait for Clk_period;
		Addr <=  "00001110111011";
		Trees_din <= x"00760f25";
		wait for Clk_period;
		Addr <=  "00001110111100";
		Trees_din <= x"03fbd804";
		wait for Clk_period;
		Addr <=  "00001110111101";
		Trees_din <= x"ffd50f25";
		wait for Clk_period;
		Addr <=  "00001110111110";
		Trees_din <= x"003b0f25";
		wait for Clk_period;
		Addr <=  "00001110111111";
		Trees_din <= x"06fc2008";
		wait for Clk_period;
		Addr <=  "00001111000000";
		Trees_din <= x"1c003804";
		wait for Clk_period;
		Addr <=  "00001111000001";
		Trees_din <= x"fff30f25";
		wait for Clk_period;
		Addr <=  "00001111000010";
		Trees_din <= x"00410f25";
		wait for Clk_period;
		Addr <=  "00001111000011";
		Trees_din <= x"000b0b08";
		wait for Clk_period;
		Addr <=  "00001111000100";
		Trees_din <= x"00e9ab04";
		wait for Clk_period;
		Addr <=  "00001111000101";
		Trees_din <= x"ffbb0f25";
		wait for Clk_period;
		Addr <=  "00001111000110";
		Trees_din <= x"00370f25";
		wait for Clk_period;
		Addr <=  "00001111000111";
		Trees_din <= x"ffa90f25";
		wait for Clk_period;
		Addr <=  "00001111001000";
		Trees_din <= x"00770f25";
		wait for Clk_period;
		Addr <=  "00001111001001";
		Trees_din <= x"050d5a28";
		wait for Clk_period;
		Addr <=  "00001111001010";
		Trees_din <= x"05039508";
		wait for Clk_period;
		Addr <=  "00001111001011";
		Trees_din <= x"0b040204";
		wait for Clk_period;
		Addr <=  "00001111001100";
		Trees_din <= x"ff800f91";
		wait for Clk_period;
		Addr <=  "00001111001101";
		Trees_din <= x"000e0f91";
		wait for Clk_period;
		Addr <=  "00001111001110";
		Trees_din <= x"09faf108";
		wait for Clk_period;
		Addr <=  "00001111001111";
		Trees_din <= x"0a01b404";
		wait for Clk_period;
		Addr <=  "00001111010000";
		Trees_din <= x"fff20f91";
		wait for Clk_period;
		Addr <=  "00001111010001";
		Trees_din <= x"00520f91";
		wait for Clk_period;
		Addr <=  "00001111010010";
		Trees_din <= x"09053410";
		wait for Clk_period;
		Addr <=  "00001111010011";
		Trees_din <= x"000b0b08";
		wait for Clk_period;
		Addr <=  "00001111010100";
		Trees_din <= x"00010e04";
		wait for Clk_period;
		Addr <=  "00001111010101";
		Trees_din <= x"ffc50f91";
		wait for Clk_period;
		Addr <=  "00001111010110";
		Trees_din <= x"00310f91";
		wait for Clk_period;
		Addr <=  "00001111010111";
		Trees_din <= x"13028604";
		wait for Clk_period;
		Addr <=  "00001111011000";
		Trees_din <= x"ff970f91";
		wait for Clk_period;
		Addr <=  "00001111011001";
		Trees_din <= x"ffe80f91";
		wait for Clk_period;
		Addr <=  "00001111011010";
		Trees_din <= x"0eff8804";
		wait for Clk_period;
		Addr <=  "00001111011011";
		Trees_din <= x"00380f91";
		wait for Clk_period;
		Addr <=  "00001111011100";
		Trees_din <= x"00060f91";
		wait for Clk_period;
		Addr <=  "00001111011101";
		Trees_din <= x"0408d30c";
		wait for Clk_period;
		Addr <=  "00001111011110";
		Trees_din <= x"000b0b04";
		wait for Clk_period;
		Addr <=  "00001111011111";
		Trees_din <= x"007b0f91";
		wait for Clk_period;
		Addr <=  "00001111100000";
		Trees_din <= x"18003804";
		wait for Clk_period;
		Addr <=  "00001111100001";
		Trees_din <= x"003c0f91";
		wait for Clk_period;
		Addr <=  "00001111100010";
		Trees_din <= x"fff30f91";
		wait for Clk_period;
		Addr <=  "00001111100011";
		Trees_din <= x"fffd0f91";
		wait for Clk_period;
		Addr <=  "00001111100100";
		Trees_din <= x"05085510";
		wait for Clk_period;
		Addr <=  "00001111100101";
		Trees_din <= x"18004e0c";
		wait for Clk_period;
		Addr <=  "00001111100110";
		Trees_din <= x"0b040208";
		wait for Clk_period;
		Addr <=  "00001111100111";
		Trees_din <= x"0506f704";
		wait for Clk_period;
		Addr <=  "00001111101000";
		Trees_din <= x"ff810ff5";
		wait for Clk_period;
		Addr <=  "00001111101001";
		Trees_din <= x"ffe60ff5";
		wait for Clk_period;
		Addr <=  "00001111101010";
		Trees_din <= x"00140ff5";
		wait for Clk_period;
		Addr <=  "00001111101011";
		Trees_din <= x"00210ff5";
		wait for Clk_period;
		Addr <=  "00001111101100";
		Trees_din <= x"05109320";
		wait for Clk_period;
		Addr <=  "00001111101101";
		Trees_din <= x"03fcf114";
		wait for Clk_period;
		Addr <=  "00001111101110";
		Trees_din <= x"08005108";
		wait for Clk_period;
		Addr <=  "00001111101111";
		Trees_din <= x"07005604";
		wait for Clk_period;
		Addr <=  "00001111110000";
		Trees_din <= x"00200ff5";
		wait for Clk_period;
		Addr <=  "00001111110001";
		Trees_din <= x"ffc70ff5";
		wait for Clk_period;
		Addr <=  "00001111110010";
		Trees_din <= x"06fcf608";
		wait for Clk_period;
		Addr <=  "00001111110011";
		Trees_din <= x"1b01aa04";
		wait for Clk_period;
		Addr <=  "00001111110100";
		Trees_din <= x"00430ff5";
		wait for Clk_period;
		Addr <=  "00001111110101";
		Trees_din <= x"fff70ff5";
		wait for Clk_period;
		Addr <=  "00001111110110";
		Trees_din <= x"00650ff5";
		wait for Clk_period;
		Addr <=  "00001111110111";
		Trees_din <= x"06fc2004";
		wait for Clk_period;
		Addr <=  "00001111111000";
		Trees_din <= x"001d0ff5";
		wait for Clk_period;
		Addr <=  "00001111111001";
		Trees_din <= x"18003b04";
		wait for Clk_period;
		Addr <=  "00001111111010";
		Trees_din <= x"fffe0ff5";
		wait for Clk_period;
		Addr <=  "00001111111011";
		Trees_din <= x"ffb50ff5";
		wait for Clk_period;
		Addr <=  "00001111111100";
		Trees_din <= x"006b0ff5";
		wait for Clk_period;
		Addr <=  "00001111111101";
		Trees_din <= x"050d5a2c";
		wait for Clk_period;
		Addr <=  "00001111111110";
		Trees_din <= x"05039508";
		wait for Clk_period;
		Addr <=  "00001111111111";
		Trees_din <= x"0f03fb04";
		wait for Clk_period;
		Addr <=  "00010000000000";
		Trees_din <= x"ff8a1061";
		wait for Clk_period;
		Addr <=  "00010000000001";
		Trees_din <= x"00101061";
		wait for Clk_period;
		Addr <=  "00010000000010";
		Trees_din <= x"1d00b10c";
		wait for Clk_period;
		Addr <=  "00010000000011";
		Trees_din <= x"03fd0f08";
		wait for Clk_period;
		Addr <=  "00010000000100";
		Trees_din <= x"07005804";
		wait for Clk_period;
		Addr <=  "00010000000101";
		Trees_din <= x"000e1061";
		wait for Clk_period;
		Addr <=  "00010000000110";
		Trees_din <= x"00531061";
		wait for Clk_period;
		Addr <=  "00010000000111";
		Trees_din <= x"fff51061";
		wait for Clk_period;
		Addr <=  "00010000001000";
		Trees_din <= x"06fdb40c";
		wait for Clk_period;
		Addr <=  "00010000001001";
		Trees_din <= x"09fad804";
		wait for Clk_period;
		Addr <=  "00010000001010";
		Trees_din <= x"000f1061";
		wait for Clk_period;
		Addr <=  "00010000001011";
		Trees_din <= x"000bb804";
		wait for Clk_period;
		Addr <=  "00010000001100";
		Trees_din <= x"ffe81061";
		wait for Clk_period;
		Addr <=  "00010000001101";
		Trees_din <= x"ff9e1061";
		wait for Clk_period;
		Addr <=  "00010000001110";
		Trees_din <= x"04ffe708";
		wait for Clk_period;
		Addr <=  "00010000001111";
		Trees_din <= x"04ff0f04";
		wait for Clk_period;
		Addr <=  "00010000010000";
		Trees_din <= x"00011061";
		wait for Clk_period;
		Addr <=  "00010000010001";
		Trees_din <= x"00461061";
		wait for Clk_period;
		Addr <=  "00010000010010";
		Trees_din <= x"ffcf1061";
		wait for Clk_period;
		Addr <=  "00010000010011";
		Trees_din <= x"0403e808";
		wait for Clk_period;
		Addr <=  "00010000010100";
		Trees_din <= x"000b0b04";
		wait for Clk_period;
		Addr <=  "00010000010101";
		Trees_din <= x"00721061";
		wait for Clk_period;
		Addr <=  "00010000010110";
		Trees_din <= x"001e1061";
		wait for Clk_period;
		Addr <=  "00010000010111";
		Trees_din <= x"00101061";
		wait for Clk_period;
		Addr <=  "00010000011000";
		Trees_din <= x"05085510";
		wait for Clk_period;
		Addr <=  "00010000011001";
		Trees_din <= x"15f97c04";
		wait for Clk_period;
		Addr <=  "00010000011010";
		Trees_din <= x"001a10bd";
		wait for Clk_period;
		Addr <=  "00010000011011";
		Trees_din <= x"0a02fb04";
		wait for Clk_period;
		Addr <=  "00010000011100";
		Trees_din <= x"ff9410bd";
		wait for Clk_period;
		Addr <=  "00010000011101";
		Trees_din <= x"1b019004";
		wait for Clk_period;
		Addr <=  "00010000011110";
		Trees_din <= x"ffda10bd";
		wait for Clk_period;
		Addr <=  "00010000011111";
		Trees_din <= x"001110bd";
		wait for Clk_period;
		Addr <=  "00010000100000";
		Trees_din <= x"0510931c";
		wait for Clk_period;
		Addr <=  "00010000100001";
		Trees_din <= x"03fcf110";
		wait for Clk_period;
		Addr <=  "00010000100010";
		Trees_din <= x"08005104";
		wait for Clk_period;
		Addr <=  "00010000100011";
		Trees_din <= x"fff210bd";
		wait for Clk_period;
		Addr <=  "00010000100100";
		Trees_din <= x"06fcf608";
		wait for Clk_period;
		Addr <=  "00010000100101";
		Trees_din <= x"000c1004";
		wait for Clk_period;
		Addr <=  "00010000100110";
		Trees_din <= x"003a10bd";
		wait for Clk_period;
		Addr <=  "00010000100111";
		Trees_din <= x"fff310bd";
		wait for Clk_period;
		Addr <=  "00010000101000";
		Trees_din <= x"005f10bd";
		wait for Clk_period;
		Addr <=  "00010000101001";
		Trees_din <= x"13028708";
		wait for Clk_period;
		Addr <=  "00010000101010";
		Trees_din <= x"13fafe04";
		wait for Clk_period;
		Addr <=  "00010000101011";
		Trees_din <= x"001210bd";
		wait for Clk_period;
		Addr <=  "00010000101100";
		Trees_din <= x"ffbf10bd";
		wait for Clk_period;
		Addr <=  "00010000101101";
		Trees_din <= x"002010bd";
		wait for Clk_period;
		Addr <=  "00010000101110";
		Trees_din <= x"006110bd";
		wait for Clk_period;
		Addr <=  "00010000101111";
		Trees_din <= x"050d5a24";
		wait for Clk_period;
		Addr <=  "00010000110000";
		Trees_din <= x"03ff7720";
		wait for Clk_period;
		Addr <=  "00010000110001";
		Trees_din <= x"1d00b108";
		wait for Clk_period;
		Addr <=  "00010000110010";
		Trees_din <= x"01fbb404";
		wait for Clk_period;
		Addr <=  "00010000110011";
		Trees_din <= x"004c1119";
		wait for Clk_period;
		Addr <=  "00010000110100";
		Trees_din <= x"fff51119";
		wait for Clk_period;
		Addr <=  "00010000110101";
		Trees_din <= x"000b6410";
		wait for Clk_period;
		Addr <=  "00010000110110";
		Trees_din <= x"0f028408";
		wait for Clk_period;
		Addr <=  "00010000110111";
		Trees_din <= x"04fe7c04";
		wait for Clk_period;
		Addr <=  "00010000111000";
		Trees_din <= x"fff81119";
		wait for Clk_period;
		Addr <=  "00010000111001";
		Trees_din <= x"ffc91119";
		wait for Clk_period;
		Addr <=  "00010000111010";
		Trees_din <= x"18003204";
		wait for Clk_period;
		Addr <=  "00010000111011";
		Trees_din <= x"00531119";
		wait for Clk_period;
		Addr <=  "00010000111100";
		Trees_din <= x"000f1119";
		wait for Clk_period;
		Addr <=  "00010000111101";
		Trees_din <= x"0f014304";
		wait for Clk_period;
		Addr <=  "00010000111110";
		Trees_din <= x"fffb1119";
		wait for Clk_period;
		Addr <=  "00010000111111";
		Trees_din <= x"ffa31119";
		wait for Clk_period;
		Addr <=  "00010001000000";
		Trees_din <= x"ffa61119";
		wait for Clk_period;
		Addr <=  "00010001000001";
		Trees_din <= x"0403e808";
		wait for Clk_period;
		Addr <=  "00010001000010";
		Trees_din <= x"000b0b04";
		wait for Clk_period;
		Addr <=  "00010001000011";
		Trees_din <= x"00681119";
		wait for Clk_period;
		Addr <=  "00010001000100";
		Trees_din <= x"001c1119";
		wait for Clk_period;
		Addr <=  "00010001000101";
		Trees_din <= x"000d1119";
		wait for Clk_period;
		Addr <=  "00010001000110";
		Trees_din <= x"0508550c";
		wait for Clk_period;
		Addr <=  "00010001000111";
		Trees_din <= x"15f97c04";
		wait for Clk_period;
		Addr <=  "00010001001000";
		Trees_din <= x"0016116d";
		wait for Clk_period;
		Addr <=  "00010001001001";
		Trees_din <= x"0a02fb04";
		wait for Clk_period;
		Addr <=  "00010001001010";
		Trees_din <= x"ff9d116d";
		wait for Clk_period;
		Addr <=  "00010001001011";
		Trees_din <= x"fff6116d";
		wait for Clk_period;
		Addr <=  "00010001001100";
		Trees_din <= x"0510931c";
		wait for Clk_period;
		Addr <=  "00010001001101";
		Trees_din <= x"0800540c";
		wait for Clk_period;
		Addr <=  "00010001001110";
		Trees_din <= x"07005608";
		wait for Clk_period;
		Addr <=  "00010001001111";
		Trees_din <= x"01fa7a04";
		wait for Clk_period;
		Addr <=  "00010001010000";
		Trees_din <= x"ffef116d";
		wait for Clk_period;
		Addr <=  "00010001010001";
		Trees_din <= x"002b116d";
		wait for Clk_period;
		Addr <=  "00010001010010";
		Trees_din <= x"ffc6116d";
		wait for Clk_period;
		Addr <=  "00010001010011";
		Trees_din <= x"1103880c";
		wait for Clk_period;
		Addr <=  "00010001010100";
		Trees_din <= x"0f028708";
		wait for Clk_period;
		Addr <=  "00010001010101";
		Trees_din <= x"04fe7c04";
		wait for Clk_period;
		Addr <=  "00010001010110";
		Trees_din <= x"005d116d";
		wait for Clk_period;
		Addr <=  "00010001010111";
		Trees_din <= x"000f116d";
		wait for Clk_period;
		Addr <=  "00010001011000";
		Trees_din <= x"0001116d";
		wait for Clk_period;
		Addr <=  "00010001011001";
		Trees_din <= x"fff4116d";
		wait for Clk_period;
		Addr <=  "00010001011010";
		Trees_din <= x"0058116d";
		wait for Clk_period;
		Addr <=  "00010001011011";
		Trees_din <= x"0506f708";
		wait for Clk_period;
		Addr <=  "00010001011100";
		Trees_din <= x"0e017f04";
		wait for Clk_period;
		Addr <=  "00010001011101";
		Trees_din <= x"ffa111b9";
		wait for Clk_period;
		Addr <=  "00010001011110";
		Trees_din <= x"001111b9";
		wait for Clk_period;
		Addr <=  "00010001011111";
		Trees_din <= x"0510931c";
		wait for Clk_period;
		Addr <=  "00010001100000";
		Trees_din <= x"03fcf110";
		wait for Clk_period;
		Addr <=  "00010001100001";
		Trees_din <= x"0a013b08";
		wait for Clk_period;
		Addr <=  "00010001100010";
		Trees_din <= x"050c4e04";
		wait for Clk_period;
		Addr <=  "00010001100011";
		Trees_din <= x"ffd211b9";
		wait for Clk_period;
		Addr <=  "00010001100100";
		Trees_din <= x"003311b9";
		wait for Clk_period;
		Addr <=  "00010001100101";
		Trees_din <= x"12009404";
		wait for Clk_period;
		Addr <=  "00010001100110";
		Trees_din <= x"006211b9";
		wait for Clk_period;
		Addr <=  "00010001100111";
		Trees_din <= x"000611b9";
		wait for Clk_period;
		Addr <=  "00010001101000";
		Trees_din <= x"06fc2004";
		wait for Clk_period;
		Addr <=  "00010001101001";
		Trees_din <= x"001911b9";
		wait for Clk_period;
		Addr <=  "00010001101010";
		Trees_din <= x"000b0b04";
		wait for Clk_period;
		Addr <=  "00010001101011";
		Trees_din <= x"fff911b9";
		wait for Clk_period;
		Addr <=  "00010001101100";
		Trees_din <= x"ffb811b9";
		wait for Clk_period;
		Addr <=  "00010001101101";
		Trees_din <= x"005211b9";
		wait for Clk_period;
		Addr <=  "00010001101110";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00010001101111";
		Trees_din <= x"0508550c";
		wait for Clk_period;
		Addr <=  "00010001110000";
		Trees_din <= x"0e017f08";
		wait for Clk_period;
		Addr <=  "00010001110001";
		Trees_din <= x"03fbcb04";
		wait for Clk_period;
		Addr <=  "00010001110010";
		Trees_din <= x"00081201";
		wait for Clk_period;
		Addr <=  "00010001110011";
		Trees_din <= x"ff9e1201";
		wait for Clk_period;
		Addr <=  "00010001110100";
		Trees_din <= x"000c1201";
		wait for Clk_period;
		Addr <=  "00010001110101";
		Trees_din <= x"05109314";
		wait for Clk_period;
		Addr <=  "00010001110110";
		Trees_din <= x"00f0ae04";
		wait for Clk_period;
		Addr <=  "00010001110111";
		Trees_din <= x"ffd21201";
		wait for Clk_period;
		Addr <=  "00010001111000";
		Trees_din <= x"08005104";
		wait for Clk_period;
		Addr <=  "00010001111001";
		Trees_din <= x"ffed1201";
		wait for Clk_period;
		Addr <=  "00010001111010";
		Trees_din <= x"0b028808";
		wait for Clk_period;
		Addr <=  "00010001111011";
		Trees_din <= x"0a02f304";
		wait for Clk_period;
		Addr <=  "00010001111100";
		Trees_din <= x"00471201";
		wait for Clk_period;
		Addr <=  "00010001111101";
		Trees_din <= x"00061201";
		wait for Clk_period;
		Addr <=  "00010001111110";
		Trees_din <= x"fff81201";
		wait for Clk_period;
		Addr <=  "00010001111111";
		Trees_din <= x"004d1201";
		wait for Clk_period;
		Addr <=  "00010010000000";
		Trees_din <= x"05039508";
		wait for Clk_period;
		Addr <=  "00010010000001";
		Trees_din <= x"0b026d04";
		wait for Clk_period;
		Addr <=  "00010010000010";
		Trees_din <= x"ffae1255";
		wait for Clk_period;
		Addr <=  "00010010000011";
		Trees_din <= x"ffef1255";
		wait for Clk_period;
		Addr <=  "00010010000100";
		Trees_din <= x"050d5a18";
		wait for Clk_period;
		Addr <=  "00010010000101";
		Trees_din <= x"0c004508";
		wait for Clk_period;
		Addr <=  "00010010000110";
		Trees_din <= x"01fae604";
		wait for Clk_period;
		Addr <=  "00010010000111";
		Trees_din <= x"00481255";
		wait for Clk_period;
		Addr <=  "00010010001000";
		Trees_din <= x"00011255";
		wait for Clk_period;
		Addr <=  "00010010001001";
		Trees_din <= x"01fa7a04";
		wait for Clk_period;
		Addr <=  "00010010001010";
		Trees_din <= x"ffc91255";
		wait for Clk_period;
		Addr <=  "00010010001011";
		Trees_din <= x"00043504";
		wait for Clk_period;
		Addr <=  "00010010001100";
		Trees_din <= x"ffd71255";
		wait for Clk_period;
		Addr <=  "00010010001101";
		Trees_din <= x"08005704";
		wait for Clk_period;
		Addr <=  "00010010001110";
		Trees_din <= x"ffff1255";
		wait for Clk_period;
		Addr <=  "00010010001111";
		Trees_din <= x"00311255";
		wait for Clk_period;
		Addr <=  "00010010010000";
		Trees_din <= x"03fcc704";
		wait for Clk_period;
		Addr <=  "00010010010001";
		Trees_din <= x"00571255";
		wait for Clk_period;
		Addr <=  "00010010010010";
		Trees_din <= x"0515e904";
		wait for Clk_period;
		Addr <=  "00010010010011";
		Trees_din <= x"ffe91255";
		wait for Clk_period;
		Addr <=  "00010010010100";
		Trees_din <= x"00401255";
		wait for Clk_period;
		Addr <=  "00010010010101";
		Trees_din <= x"05039504";
		wait for Clk_period;
		Addr <=  "00010010010110";
		Trees_din <= x"ffc212a1";
		wait for Clk_period;
		Addr <=  "00010010010111";
		Trees_din <= x"050d5a18";
		wait for Clk_period;
		Addr <=  "00010010011000";
		Trees_din <= x"0c00910c";
		wait for Clk_period;
		Addr <=  "00010010011001";
		Trees_din <= x"0f00bc04";
		wait for Clk_period;
		Addr <=  "00010010011010";
		Trees_din <= x"ffec12a1";
		wait for Clk_period;
		Addr <=  "00010010011011";
		Trees_din <= x"01fbd304";
		wait for Clk_period;
		Addr <=  "00010010011100";
		Trees_din <= x"003f12a1";
		wait for Clk_period;
		Addr <=  "00010010011101";
		Trees_din <= x"000f12a1";
		wait for Clk_period;
		Addr <=  "00010010011110";
		Trees_din <= x"06fdf108";
		wait for Clk_period;
		Addr <=  "00010010011111";
		Trees_din <= x"04fe2204";
		wait for Clk_period;
		Addr <=  "00010010100000";
		Trees_din <= x"000212a1";
		wait for Clk_period;
		Addr <=  "00010010100001";
		Trees_din <= x"ffb512a1";
		wait for Clk_period;
		Addr <=  "00010010100010";
		Trees_din <= x"000812a1";
		wait for Clk_period;
		Addr <=  "00010010100011";
		Trees_din <= x"0403e808";
		wait for Clk_period;
		Addr <=  "00010010100100";
		Trees_din <= x"000b0b04";
		wait for Clk_period;
		Addr <=  "00010010100101";
		Trees_din <= x"005712a1";
		wait for Clk_period;
		Addr <=  "00010010100110";
		Trees_din <= x"001612a1";
		wait for Clk_period;
		Addr <=  "00010010100111";
		Trees_din <= x"000412a1";
		wait for Clk_period;
		Addr <=  "00010010101000";
		Trees_din <= x"0508550c";
		wait for Clk_period;
		Addr <=  "00010010101001";
		Trees_din <= x"0e017f08";
		wait for Clk_period;
		Addr <=  "00010010101010";
		Trees_din <= x"03fc0304";
		wait for Clk_period;
		Addr <=  "00010010101011";
		Trees_din <= x"000312ed";
		wait for Clk_period;
		Addr <=  "00010010101100";
		Trees_din <= x"ffaa12ed";
		wait for Clk_period;
		Addr <=  "00010010101101";
		Trees_din <= x"000e12ed";
		wait for Clk_period;
		Addr <=  "00010010101110";
		Trees_din <= x"05109318";
		wait for Clk_period;
		Addr <=  "00010010101111";
		Trees_din <= x"03fcf10c";
		wait for Clk_period;
		Addr <=  "00010010110000";
		Trees_din <= x"0a008604";
		wait for Clk_period;
		Addr <=  "00010010110001";
		Trees_din <= x"fff112ed";
		wait for Clk_period;
		Addr <=  "00010010110010";
		Trees_din <= x"0f007904";
		wait for Clk_period;
		Addr <=  "00010010110011";
		Trees_din <= x"000e12ed";
		wait for Clk_period;
		Addr <=  "00010010110100";
		Trees_din <= x"004512ed";
		wait for Clk_period;
		Addr <=  "00010010110101";
		Trees_din <= x"06fc2004";
		wait for Clk_period;
		Addr <=  "00010010110110";
		Trees_din <= x"001312ed";
		wait for Clk_period;
		Addr <=  "00010010110111";
		Trees_din <= x"18003b04";
		wait for Clk_period;
		Addr <=  "00010010111000";
		Trees_din <= x"000012ed";
		wait for Clk_period;
		Addr <=  "00010010111001";
		Trees_din <= x"ffc312ed";
		wait for Clk_period;
		Addr <=  "00010010111010";
		Trees_din <= x"004312ed";
		wait for Clk_period;
		Addr <=  "00010010111011";
		Trees_din <= x"05072408";
		wait for Clk_period;
		Addr <=  "00010010111100";
		Trees_din <= x"0f037904";
		wait for Clk_period;
		Addr <=  "00010010111101";
		Trees_din <= x"ffba1331";
		wait for Clk_period;
		Addr <=  "00010010111110";
		Trees_din <= x"000d1331";
		wait for Clk_period;
		Addr <=  "00010010111111";
		Trees_din <= x"03fcf110";
		wait for Clk_period;
		Addr <=  "00010011000000";
		Trees_din <= x"0a013b08";
		wait for Clk_period;
		Addr <=  "00010011000001";
		Trees_din <= x"050c4e04";
		wait for Clk_period;
		Addr <=  "00010011000010";
		Trees_din <= x"ffd81331";
		wait for Clk_period;
		Addr <=  "00010011000011";
		Trees_din <= x"00371331";
		wait for Clk_period;
		Addr <=  "00010011000100";
		Trees_din <= x"12009404";
		wait for Clk_period;
		Addr <=  "00010011000101";
		Trees_din <= x"00581331";
		wait for Clk_period;
		Addr <=  "00010011000110";
		Trees_din <= x"00101331";
		wait for Clk_period;
		Addr <=  "00010011000111";
		Trees_din <= x"000b0b08";
		wait for Clk_period;
		Addr <=  "00010011001000";
		Trees_din <= x"04086d04";
		wait for Clk_period;
		Addr <=  "00010011001001";
		Trees_din <= x"00351331";
		wait for Clk_period;
		Addr <=  "00010011001010";
		Trees_din <= x"ffe71331";
		wait for Clk_period;
		Addr <=  "00010011001011";
		Trees_din <= x"ffdd1331";
		wait for Clk_period;
		Addr <=  "00010011001100";
		Trees_din <= x"050d5a18";
		wait for Clk_period;
		Addr <=  "00010011001101";
		Trees_din <= x"01027c14";
		wait for Clk_period;
		Addr <=  "00010011001110";
		Trees_din <= x"000b6408";
		wait for Clk_period;
		Addr <=  "00010011001111";
		Trees_din <= x"0f028704";
		wait for Clk_period;
		Addr <=  "00010011010000";
		Trees_din <= x"fff61375";
		wait for Clk_period;
		Addr <=  "00010011010001";
		Trees_din <= x"00451375";
		wait for Clk_period;
		Addr <=  "00010011010010";
		Trees_din <= x"09fa5304";
		wait for Clk_period;
		Addr <=  "00010011010011";
		Trees_din <= x"00241375";
		wait for Clk_period;
		Addr <=  "00010011010100";
		Trees_din <= x"0904ba04";
		wait for Clk_period;
		Addr <=  "00010011010101";
		Trees_din <= x"ffaa1375";
		wait for Clk_period;
		Addr <=  "00010011010110";
		Trees_din <= x"000d1375";
		wait for Clk_period;
		Addr <=  "00010011010111";
		Trees_din <= x"ffb71375";
		wait for Clk_period;
		Addr <=  "00010011011000";
		Trees_din <= x"0d011b04";
		wait for Clk_period;
		Addr <=  "00010011011001";
		Trees_din <= x"00081375";
		wait for Clk_period;
		Addr <=  "00010011011010";
		Trees_din <= x"15028604";
		wait for Clk_period;
		Addr <=  "00010011011011";
		Trees_din <= x"00151375";
		wait for Clk_period;
		Addr <=  "00010011011100";
		Trees_din <= x"00511375";
		wait for Clk_period;
		Addr <=  "00010011011101";
		Trees_din <= x"050d5a18";
		wait for Clk_period;
		Addr <=  "00010011011110";
		Trees_din <= x"01007714";
		wait for Clk_period;
		Addr <=  "00010011011111";
		Trees_din <= x"1000a704";
		wait for Clk_period;
		Addr <=  "00010011100000";
		Trees_din <= x"ffdb13b9";
		wait for Clk_period;
		Addr <=  "00010011100001";
		Trees_din <= x"02fd8604";
		wait for Clk_period;
		Addr <=  "00010011100010";
		Trees_din <= x"ffe213b9";
		wait for Clk_period;
		Addr <=  "00010011100011";
		Trees_din <= x"000b0b04";
		wait for Clk_period;
		Addr <=  "00010011100100";
		Trees_din <= x"004013b9";
		wait for Clk_period;
		Addr <=  "00010011100101";
		Trees_din <= x"1b026804";
		wait for Clk_period;
		Addr <=  "00010011100110";
		Trees_din <= x"ffe613b9";
		wait for Clk_period;
		Addr <=  "00010011100111";
		Trees_din <= x"002313b9";
		wait for Clk_period;
		Addr <=  "00010011101000";
		Trees_din <= x"ffbf13b9";
		wait for Clk_period;
		Addr <=  "00010011101001";
		Trees_din <= x"0403e808";
		wait for Clk_period;
		Addr <=  "00010011101010";
		Trees_din <= x"000b0b04";
		wait for Clk_period;
		Addr <=  "00010011101011";
		Trees_din <= x"004b13b9";
		wait for Clk_period;
		Addr <=  "00010011101100";
		Trees_din <= x"001613b9";
		wait for Clk_period;
		Addr <=  "00010011101101";
		Trees_din <= x"000413b9";
		wait for Clk_period;
		Addr <=  "00010011101110";
		Trees_din <= x"0508550c";
		wait for Clk_period;
		Addr <=  "00010011101111";
		Trees_din <= x"0e017f08";
		wait for Clk_period;
		Addr <=  "00010011110000";
		Trees_din <= x"17004504";
		wait for Clk_period;
		Addr <=  "00010011110001";
		Trees_din <= x"ffb713f5";
		wait for Clk_period;
		Addr <=  "00010011110010";
		Trees_din <= x"fff913f5";
		wait for Clk_period;
		Addr <=  "00010011110011";
		Trees_din <= x"000713f5";
		wait for Clk_period;
		Addr <=  "00010011110100";
		Trees_din <= x"03fcf10c";
		wait for Clk_period;
		Addr <=  "00010011110101";
		Trees_din <= x"08005104";
		wait for Clk_period;
		Addr <=  "00010011110110";
		Trees_din <= x"fffb13f5";
		wait for Clk_period;
		Addr <=  "00010011110111";
		Trees_din <= x"0f007904";
		wait for Clk_period;
		Addr <=  "00010011111000";
		Trees_din <= x"001313f5";
		wait for Clk_period;
		Addr <=  "00010011111001";
		Trees_din <= x"004b13f5";
		wait for Clk_period;
		Addr <=  "00010011111010";
		Trees_din <= x"00087604";
		wait for Clk_period;
		Addr <=  "00010011111011";
		Trees_din <= x"001a13f5";
		wait for Clk_period;
		Addr <=  "00010011111100";
		Trees_din <= x"ffe913f5";
		wait for Clk_period;
		Addr <=  "00010011111101";
		Trees_din <= x"0507e108";
		wait for Clk_period;
		Addr <=  "00010011111110";
		Trees_din <= x"10028704";
		wait for Clk_period;
		Addr <=  "00010011111111";
		Trees_din <= x"ffc81429";
		wait for Clk_period;
		Addr <=  "00010100000000";
		Trees_din <= x"00021429";
		wait for Clk_period;
		Addr <=  "00010100000001";
		Trees_din <= x"050d5a0c";
		wait for Clk_period;
		Addr <=  "00010100000010";
		Trees_din <= x"08005404";
		wait for Clk_period;
		Addr <=  "00010100000011";
		Trees_din <= x"ffe31429";
		wait for Clk_period;
		Addr <=  "00010100000100";
		Trees_din <= x"0d01b604";
		wait for Clk_period;
		Addr <=  "00010100000101";
		Trees_din <= x"fffc1429";
		wait for Clk_period;
		Addr <=  "00010100000110";
		Trees_din <= x"00301429";
		wait for Clk_period;
		Addr <=  "00010100000111";
		Trees_din <= x"0d011b04";
		wait for Clk_period;
		Addr <=  "00010100001000";
		Trees_din <= x"00061429";
		wait for Clk_period;
		Addr <=  "00010100001001";
		Trees_din <= x"003f1429";
		wait for Clk_period;
		Addr <=  "00010100001010";
		Trees_din <= x"0506f708";
		wait for Clk_period;
		Addr <=  "00010100001011";
		Trees_din <= x"0f02b804";
		wait for Clk_period;
		Addr <=  "00010100001100";
		Trees_din <= x"ffc31465";
		wait for Clk_period;
		Addr <=  "00010100001101";
		Trees_din <= x"00011465";
		wait for Clk_period;
		Addr <=  "00010100001110";
		Trees_din <= x"03fcf10c";
		wait for Clk_period;
		Addr <=  "00010100001111";
		Trees_din <= x"0a008604";
		wait for Clk_period;
		Addr <=  "00010100010000";
		Trees_din <= x"fffc1465";
		wait for Clk_period;
		Addr <=  "00010100010001";
		Trees_din <= x"17004404";
		wait for Clk_period;
		Addr <=  "00010100010010";
		Trees_din <= x"00151465";
		wait for Clk_period;
		Addr <=  "00010100010011";
		Trees_din <= x"00451465";
		wait for Clk_period;
		Addr <=  "00010100010100";
		Trees_din <= x"0bfe7e04";
		wait for Clk_period;
		Addr <=  "00010100010101";
		Trees_din <= x"ffdd1465";
		wait for Clk_period;
		Addr <=  "00010100010110";
		Trees_din <= x"03fe4204";
		wait for Clk_period;
		Addr <=  "00010100010111";
		Trees_din <= x"fff11465";
		wait for Clk_period;
		Addr <=  "00010100011000";
		Trees_din <= x"00231465";
		wait for Clk_period;
		Addr <=  "00010100011001";
		Trees_din <= x"050d5a14";
		wait for Clk_period;
		Addr <=  "00010100011010";
		Trees_din <= x"0c004408";
		wait for Clk_period;
		Addr <=  "00010100011011";
		Trees_din <= x"1503cc04";
		wait for Clk_period;
		Addr <=  "00010100011100";
		Trees_din <= x"00031499";
		wait for Clk_period;
		Addr <=  "00010100011101";
		Trees_din <= x"00221499";
		wait for Clk_period;
		Addr <=  "00010100011110";
		Trees_din <= x"0c027008";
		wait for Clk_period;
		Addr <=  "00010100011111";
		Trees_din <= x"08005704";
		wait for Clk_period;
		Addr <=  "00010100100000";
		Trees_din <= x"ffc41499";
		wait for Clk_period;
		Addr <=  "00010100100001";
		Trees_din <= x"fffc1499";
		wait for Clk_period;
		Addr <=  "00010100100010";
		Trees_din <= x"00091499";
		wait for Clk_period;
		Addr <=  "00010100100011";
		Trees_din <= x"0d011b04";
		wait for Clk_period;
		Addr <=  "00010100100100";
		Trees_din <= x"00061499";
		wait for Clk_period;
		Addr <=  "00010100100101";
		Trees_din <= x"003c1499";
		wait for Clk_period;
		Addr <=  "00010100100110";
		Trees_din <= x"05085508";
		wait for Clk_period;
		Addr <=  "00010100100111";
		Trees_din <= x"06ff1b04";
		wait for Clk_period;
		Addr <=  "00010100101000";
		Trees_din <= x"ffcb14c5";
		wait for Clk_period;
		Addr <=  "00010100101001";
		Trees_din <= x"ffff14c5";
		wait for Clk_period;
		Addr <=  "00010100101010";
		Trees_din <= x"0b02880c";
		wait for Clk_period;
		Addr <=  "00010100101011";
		Trees_din <= x"11013104";
		wait for Clk_period;
		Addr <=  "00010100101100";
		Trees_din <= x"fffe14c5";
		wait for Clk_period;
		Addr <=  "00010100101101";
		Trees_din <= x"18003c04";
		wait for Clk_period;
		Addr <=  "00010100101110";
		Trees_din <= x"004114c5";
		wait for Clk_period;
		Addr <=  "00010100101111";
		Trees_din <= x"000a14c5";
		wait for Clk_period;
		Addr <=  "00010100110000";
		Trees_din <= x"fff514c5";
		wait for Clk_period;
		Addr <=  "00010100110001";
		Trees_din <= x"050d5a14";
		wait for Clk_period;
		Addr <=  "00010100110010";
		Trees_din <= x"01007710";
		wait for Clk_period;
		Addr <=  "00010100110011";
		Trees_din <= x"01fa2a04";
		wait for Clk_period;
		Addr <=  "00010100110100";
		Trees_din <= x"ffdf14f9";
		wait for Clk_period;
		Addr <=  "00010100110101";
		Trees_din <= x"000b6404";
		wait for Clk_period;
		Addr <=  "00010100110110";
		Trees_din <= x"002c14f9";
		wait for Clk_period;
		Addr <=  "00010100110111";
		Trees_din <= x"1b021f04";
		wait for Clk_period;
		Addr <=  "00010100111000";
		Trees_din <= x"ffea14f9";
		wait for Clk_period;
		Addr <=  "00010100111001";
		Trees_din <= x"000d14f9";
		wait for Clk_period;
		Addr <=  "00010100111010";
		Trees_din <= x"ffc514f9";
		wait for Clk_period;
		Addr <=  "00010100111011";
		Trees_din <= x"18003b04";
		wait for Clk_period;
		Addr <=  "00010100111100";
		Trees_din <= x"003714f9";
		wait for Clk_period;
		Addr <=  "00010100111101";
		Trees_din <= x"000514f9";
		wait for Clk_period;
		Addr <=  "00010100111110";
		Trees_din <= x"05072408";
		wait for Clk_period;
		Addr <=  "00010100111111";
		Trees_din <= x"16006604";
		wait for Clk_period;
		Addr <=  "00010101000000";
		Trees_din <= x"ffcf1535";
		wait for Clk_period;
		Addr <=  "00010101000001";
		Trees_din <= x"fffb1535";
		wait for Clk_period;
		Addr <=  "00010101000010";
		Trees_din <= x"03fcf10c";
		wait for Clk_period;
		Addr <=  "00010101000011";
		Trees_din <= x"08005104";
		wait for Clk_period;
		Addr <=  "00010101000100";
		Trees_din <= x"fffe1535";
		wait for Clk_period;
		Addr <=  "00010101000101";
		Trees_din <= x"06fcf604";
		wait for Clk_period;
		Addr <=  "00010101000110";
		Trees_din <= x"00121535";
		wait for Clk_period;
		Addr <=  "00010101000111";
		Trees_din <= x"003f1535";
		wait for Clk_period;
		Addr <=  "00010101001000";
		Trees_din <= x"12009204";
		wait for Clk_period;
		Addr <=  "00010101001001";
		Trees_din <= x"ffe31535";
		wait for Clk_period;
		Addr <=  "00010101001010";
		Trees_din <= x"0d01c004";
		wait for Clk_period;
		Addr <=  "00010101001011";
		Trees_din <= x"fff61535";
		wait for Clk_period;
		Addr <=  "00010101001100";
		Trees_din <= x"00231535";
		wait for Clk_period;
		Addr <=  "00010101001101";
		Trees_din <= x"050d5a10";
		wait for Clk_period;
		Addr <=  "00010101001110";
		Trees_din <= x"0c004404";
		wait for Clk_period;
		Addr <=  "00010101001111";
		Trees_din <= x"00171561";
		wait for Clk_period;
		Addr <=  "00010101010000";
		Trees_din <= x"0a013b04";
		wait for Clk_period;
		Addr <=  "00010101010001";
		Trees_din <= x"ffc91561";
		wait for Clk_period;
		Addr <=  "00010101010010";
		Trees_din <= x"16001504";
		wait for Clk_period;
		Addr <=  "00010101010011";
		Trees_din <= x"ffe41561";
		wait for Clk_period;
		Addr <=  "00010101010100";
		Trees_din <= x"001b1561";
		wait for Clk_period;
		Addr <=  "00010101010101";
		Trees_din <= x"0d011b04";
		wait for Clk_period;
		Addr <=  "00010101010110";
		Trees_din <= x"00041561";
		wait for Clk_period;
		Addr <=  "00010101010111";
		Trees_din <= x"00351561";
		wait for Clk_period;
		Addr <=  "00010101011000";
		Trees_din <= x"05085508";
		wait for Clk_period;
		Addr <=  "00010101011001";
		Trees_din <= x"06ff1b04";
		wait for Clk_period;
		Addr <=  "00010101011010";
		Trees_din <= x"ffcf1595";
		wait for Clk_period;
		Addr <=  "00010101011011";
		Trees_din <= x"fffe1595";
		wait for Clk_period;
		Addr <=  "00010101011100";
		Trees_din <= x"09fade04";
		wait for Clk_period;
		Addr <=  "00010101011101";
		Trees_din <= x"002f1595";
		wait for Clk_period;
		Addr <=  "00010101011110";
		Trees_din <= x"050d5a08";
		wait for Clk_period;
		Addr <=  "00010101011111";
		Trees_din <= x"11018404";
		wait for Clk_period;
		Addr <=  "00010101100000";
		Trees_din <= x"ffde1595";
		wait for Clk_period;
		Addr <=  "00010101100001";
		Trees_din <= x"00091595";
		wait for Clk_period;
		Addr <=  "00010101100010";
		Trees_din <= x"04ff3604";
		wait for Clk_period;
		Addr <=  "00010101100011";
		Trees_din <= x"002c1595";
		wait for Clk_period;
		Addr <=  "00010101100100";
		Trees_din <= x"ffff1595";
		wait for Clk_period;
		Addr <=  "00010101100101";
		Trees_din <= x"05039504";
		wait for Clk_period;
		Addr <=  "00010101100110";
		Trees_din <= x"ffd315c9";
		wait for Clk_period;
		Addr <=  "00010101100111";
		Trees_din <= x"0c017510";
		wait for Clk_period;
		Addr <=  "00010101101000";
		Trees_din <= x"04002a0c";
		wait for Clk_period;
		Addr <=  "00010101101001";
		Trees_din <= x"000b0b04";
		wait for Clk_period;
		Addr <=  "00010101101010";
		Trees_din <= x"004515c9";
		wait for Clk_period;
		Addr <=  "00010101101011";
		Trees_din <= x"15042d04";
		wait for Clk_period;
		Addr <=  "00010101101100";
		Trees_din <= x"fff815c9";
		wait for Clk_period;
		Addr <=  "00010101101101";
		Trees_din <= x"002415c9";
		wait for Clk_period;
		Addr <=  "00010101101110";
		Trees_din <= x"ffeb15c9";
		wait for Clk_period;
		Addr <=  "00010101101111";
		Trees_din <= x"1d00e304";
		wait for Clk_period;
		Addr <=  "00010101110000";
		Trees_din <= x"ffda15c9";
		wait for Clk_period;
		Addr <=  "00010101110001";
		Trees_din <= x"001615c9";
		wait for Clk_period;
		Addr <=  "00010101110010";
		Trees_din <= x"05085508";
		wait for Clk_period;
		Addr <=  "00010101110011";
		Trees_din <= x"0f028704";
		wait for Clk_period;
		Addr <=  "00010101110100";
		Trees_din <= x"ffd315f5";
		wait for Clk_period;
		Addr <=  "00010101110101";
		Trees_din <= x"000115f5";
		wait for Clk_period;
		Addr <=  "00010101110110";
		Trees_din <= x"03fcf108";
		wait for Clk_period;
		Addr <=  "00010101110111";
		Trees_din <= x"08005304";
		wait for Clk_period;
		Addr <=  "00010101111000";
		Trees_din <= x"000315f5";
		wait for Clk_period;
		Addr <=  "00010101111001";
		Trees_din <= x"003215f5";
		wait for Clk_period;
		Addr <=  "00010101111010";
		Trees_din <= x"000b0b04";
		wait for Clk_period;
		Addr <=  "00010101111011";
		Trees_din <= x"001015f5";
		wait for Clk_period;
		Addr <=  "00010101111100";
		Trees_din <= x"ffe915f5";
		wait for Clk_period;
		Addr <=  "00010101111101";
		Trees_din <= x"05072404";
		wait for Clk_period;
		Addr <=  "00010101111110";
		Trees_din <= x"ffe01619";
		wait for Clk_period;
		Addr <=  "00010101111111";
		Trees_din <= x"04fe7c08";
		wait for Clk_period;
		Addr <=  "00010110000000";
		Trees_din <= x"08005204";
		wait for Clk_period;
		Addr <=  "00010110000001";
		Trees_din <= x"fff41619";
		wait for Clk_period;
		Addr <=  "00010110000010";
		Trees_din <= x"00311619";
		wait for Clk_period;
		Addr <=  "00010110000011";
		Trees_din <= x"1900a204";
		wait for Clk_period;
		Addr <=  "00010110000100";
		Trees_din <= x"ffe81619";
		wait for Clk_period;
		Addr <=  "00010110000101";
		Trees_din <= x"00181619";
		wait for Clk_period;
		Addr <=  "00010110000110";
		Trees_din <= x"05085508";
		wait for Clk_period;
		Addr <=  "00010110000111";
		Trees_din <= x"0f028704";
		wait for Clk_period;
		Addr <=  "00010110001000";
		Trees_din <= x"ffd61645";
		wait for Clk_period;
		Addr <=  "00010110001001";
		Trees_din <= x"00021645";
		wait for Clk_period;
		Addr <=  "00010110001010";
		Trees_din <= x"09fade04";
		wait for Clk_period;
		Addr <=  "00010110001011";
		Trees_din <= x"00291645";
		wait for Clk_period;
		Addr <=  "00010110001100";
		Trees_din <= x"050d5a08";
		wait for Clk_period;
		Addr <=  "00010110001101";
		Trees_din <= x"01fa2a04";
		wait for Clk_period;
		Addr <=  "00010110001110";
		Trees_din <= x"ffdb1645";
		wait for Clk_period;
		Addr <=  "00010110001111";
		Trees_din <= x"00021645";
		wait for Clk_period;
		Addr <=  "00010110010000";
		Trees_din <= x"001a1645";
		wait for Clk_period;
		Addr <=  "00010110010001";
		Trees_din <= x"0506f704";
		wait for Clk_period;
		Addr <=  "00010110010010";
		Trees_din <= x"ffe11671";
		wait for Clk_period;
		Addr <=  "00010110010011";
		Trees_din <= x"0b028810";
		wait for Clk_period;
		Addr <=  "00010110010100";
		Trees_din <= x"1c003208";
		wait for Clk_period;
		Addr <=  "00010110010101";
		Trees_din <= x"11013104";
		wait for Clk_period;
		Addr <=  "00010110010110";
		Trees_din <= x"ffe01671";
		wait for Clk_period;
		Addr <=  "00010110010111";
		Trees_din <= x"00191671";
		wait for Clk_period;
		Addr <=  "00010110011000";
		Trees_din <= x"03fc6b04";
		wait for Clk_period;
		Addr <=  "00010110011001";
		Trees_din <= x"003c1671";
		wait for Clk_period;
		Addr <=  "00010110011010";
		Trees_din <= x"00091671";
		wait for Clk_period;
		Addr <=  "00010110011011";
		Trees_din <= x"ffef1671";
		wait for Clk_period;
		Addr <=  "00010110011100";
		Trees_din <= x"05085508";
		wait for Clk_period;
		Addr <=  "00010110011101";
		Trees_din <= x"0f028704";
		wait for Clk_period;
		Addr <=  "00010110011110";
		Trees_din <= x"ffd9169d";
		wait for Clk_period;
		Addr <=  "00010110011111";
		Trees_din <= x"0001169d";
		wait for Clk_period;
		Addr <=  "00010110100000";
		Trees_din <= x"09fade04";
		wait for Clk_period;
		Addr <=  "00010110100001";
		Trees_din <= x"0025169d";
		wait for Clk_period;
		Addr <=  "00010110100010";
		Trees_din <= x"050d5a08";
		wait for Clk_period;
		Addr <=  "00010110100011";
		Trees_din <= x"000bb804";
		wait for Clk_period;
		Addr <=  "00010110100100";
		Trees_din <= x"0003169d";
		wait for Clk_period;
		Addr <=  "00010110100101";
		Trees_din <= x"ffde169d";
		wait for Clk_period;
		Addr <=  "00010110100110";
		Trees_din <= x"0019169d";
		wait for Clk_period;
		Addr <=  "00010110100111";
		Trees_din <= x"0c004508";
		wait for Clk_period;
		Addr <=  "00010110101000";
		Trees_din <= x"01fae604";
		wait for Clk_period;
		Addr <=  "00010110101001";
		Trees_din <= x"002d16c1";
		wait for Clk_period;
		Addr <=  "00010110101010";
		Trees_din <= x"ffff16c1";
		wait for Clk_period;
		Addr <=  "00010110101011";
		Trees_din <= x"18003908";
		wait for Clk_period;
		Addr <=  "00010110101100";
		Trees_din <= x"11013604";
		wait for Clk_period;
		Addr <=  "00010110101101";
		Trees_din <= x"ffed16c1";
		wait for Clk_period;
		Addr <=  "00010110101110";
		Trees_din <= x"001c16c1";
		wait for Clk_period;
		Addr <=  "00010110101111";
		Trees_din <= x"ffdd16c1";
		wait for Clk_period;
		Addr <=  "00010110110000";
		Trees_din <= x"05072404";
		wait for Clk_period;
		Addr <=  "00010110110001";
		Trees_din <= x"ffe516e5";
		wait for Clk_period;
		Addr <=  "00010110110010";
		Trees_din <= x"03fcf108";
		wait for Clk_period;
		Addr <=  "00010110110011";
		Trees_din <= x"0a013b04";
		wait for Clk_period;
		Addr <=  "00010110110100";
		Trees_din <= x"000216e5";
		wait for Clk_period;
		Addr <=  "00010110110101";
		Trees_din <= x"002d16e5";
		wait for Clk_period;
		Addr <=  "00010110110110";
		Trees_din <= x"12009404";
		wait for Clk_period;
		Addr <=  "00010110110111";
		Trees_din <= x"ffe616e5";
		wait for Clk_period;
		Addr <=  "00010110111000";
		Trees_din <= x"000b16e5";
		wait for Clk_period;
		Addr <=  "00010110111001";
		Trees_din <= x"0c004508";
		wait for Clk_period;
		Addr <=  "00010110111010";
		Trees_din <= x"01fae604";
		wait for Clk_period;
		Addr <=  "00010110111011";
		Trees_din <= x"002a1709";
		wait for Clk_period;
		Addr <=  "00010110111100";
		Trees_din <= x"00001709";
		wait for Clk_period;
		Addr <=  "00010110111101";
		Trees_din <= x"18003908";
		wait for Clk_period;
		Addr <=  "00010110111110";
		Trees_din <= x"1200a004";
		wait for Clk_period;
		Addr <=  "00010110111111";
		Trees_din <= x"001a1709";
		wait for Clk_period;
		Addr <=  "00010111000000";
		Trees_din <= x"ffee1709";
		wait for Clk_period;
		Addr <=  "00010111000001";
		Trees_din <= x"ffe01709";
		wait for Clk_period;
		Addr <=  "00010111000010";
		Trees_din <= x"05085504";
		wait for Clk_period;
		Addr <=  "00010111000011";
		Trees_din <= x"ffe7172d";
		wait for Clk_period;
		Addr <=  "00010111000100";
		Trees_din <= x"03fcf108";
		wait for Clk_period;
		Addr <=  "00010111000101";
		Trees_din <= x"08005304";
		wait for Clk_period;
		Addr <=  "00010111000110";
		Trees_din <= x"0000172d";
		wait for Clk_period;
		Addr <=  "00010111000111";
		Trees_din <= x"002d172d";
		wait for Clk_period;
		Addr <=  "00010111001000";
		Trees_din <= x"00087604";
		wait for Clk_period;
		Addr <=  "00010111001001";
		Trees_din <= x"000e172d";
		wait for Clk_period;
		Addr <=  "00010111001010";
		Trees_din <= x"ffec172d";
		wait for Clk_period;
		Addr <=  "00010111001011";
		Trees_din <= x"05085504";
		wait for Clk_period;
		Addr <=  "00010111001100";
		Trees_din <= x"ffe91751";
		wait for Clk_period;
		Addr <=  "00010111001101";
		Trees_din <= x"03fcf108";
		wait for Clk_period;
		Addr <=  "00010111001110";
		Trees_din <= x"08005304";
		wait for Clk_period;
		Addr <=  "00010111001111";
		Trees_din <= x"00011751";
		wait for Clk_period;
		Addr <=  "00010111010000";
		Trees_din <= x"002a1751";
		wait for Clk_period;
		Addr <=  "00010111010001";
		Trees_din <= x"03fe4204";
		wait for Clk_period;
		Addr <=  "00010111010010";
		Trees_din <= x"ffed1751";
		wait for Clk_period;
		Addr <=  "00010111010011";
		Trees_din <= x"000d1751";
		wait for Clk_period;
		Addr <=  "00010111010100";
		Trees_din <= x"01027c10";
		wait for Clk_period;
		Addr <=  "00010111010101";
		Trees_din <= x"08005204";
		wait for Clk_period;
		Addr <=  "00010111010110";
		Trees_din <= x"fff21775";
		wait for Clk_period;
		Addr <=  "00010111010111";
		Trees_din <= x"02fdf404";
		wait for Clk_period;
		Addr <=  "00010111011000";
		Trees_din <= x"fff71775";
		wait for Clk_period;
		Addr <=  "00010111011001";
		Trees_din <= x"13021e04";
		wait for Clk_period;
		Addr <=  "00010111011010";
		Trees_din <= x"002e1775";
		wait for Clk_period;
		Addr <=  "00010111011011";
		Trees_din <= x"000b1775";
		wait for Clk_period;
		Addr <=  "00010111011100";
		Trees_din <= x"ffe71775";
		wait for Clk_period;
		Addr <=  "00010111011101";
		Trees_din <= x"050d5a10";
		wait for Clk_period;
		Addr <=  "00010111011110";
		Trees_din <= x"1d00b104";
		wait for Clk_period;
		Addr <=  "00010111011111";
		Trees_din <= x"001517a1";
		wait for Clk_period;
		Addr <=  "00010111100000";
		Trees_din <= x"0f028708";
		wait for Clk_period;
		Addr <=  "00010111100001";
		Trees_din <= x"0509dd04";
		wait for Clk_period;
		Addr <=  "00010111100010";
		Trees_din <= x"ffc417a1";
		wait for Clk_period;
		Addr <=  "00010111100011";
		Trees_din <= x"fffd17a1";
		wait for Clk_period;
		Addr <=  "00010111100100";
		Trees_din <= x"000517a1";
		wait for Clk_period;
		Addr <=  "00010111100101";
		Trees_din <= x"0efe6b04";
		wait for Clk_period;
		Addr <=  "00010111100110";
		Trees_din <= x"002a17a1";
		wait for Clk_period;
		Addr <=  "00010111100111";
		Trees_din <= x"000817a1";
		wait for Clk_period;
		Addr <=  "00010111101000";
		Trees_din <= x"05072404";
		wait for Clk_period;
		Addr <=  "00010111101001";
		Trees_din <= x"ffe717c5";
		wait for Clk_period;
		Addr <=  "00010111101010";
		Trees_din <= x"04fe7c08";
		wait for Clk_period;
		Addr <=  "00010111101011";
		Trees_din <= x"08005404";
		wait for Clk_period;
		Addr <=  "00010111101100";
		Trees_din <= x"000017c5";
		wait for Clk_period;
		Addr <=  "00010111101101";
		Trees_din <= x"002b17c5";
		wait for Clk_period;
		Addr <=  "00010111101110";
		Trees_din <= x"0c008f04";
		wait for Clk_period;
		Addr <=  "00010111101111";
		Trees_din <= x"001117c5";
		wait for Clk_period;
		Addr <=  "00010111110000";
		Trees_din <= x"ffe917c5";
		wait for Clk_period;
		Addr <=  "00010111110001";
		Trees_din <= x"05085504";
		wait for Clk_period;
		Addr <=  "00010111110010";
		Trees_din <= x"ffeb17e9";
		wait for Clk_period;
		Addr <=  "00010111110011";
		Trees_din <= x"09fade04";
		wait for Clk_period;
		Addr <=  "00010111110100";
		Trees_din <= x"002217e9";
		wait for Clk_period;
		Addr <=  "00010111110101";
		Trees_din <= x"0904c908";
		wait for Clk_period;
		Addr <=  "00010111110110";
		Trees_din <= x"000b0b04";
		wait for Clk_period;
		Addr <=  "00010111110111";
		Trees_din <= x"000a17e9";
		wait for Clk_period;
		Addr <=  "00010111111000";
		Trees_din <= x"ffdc17e9";
		wait for Clk_period;
		Addr <=  "00010111111001";
		Trees_din <= x"001617e9";
		wait for Clk_period;
		Addr <=  "00010111111010";
		Trees_din <= x"04030b10";
		wait for Clk_period;
		Addr <=  "00010111111011";
		Trees_din <= x"050d5a0c";
		wait for Clk_period;
		Addr <=  "00010111111100";
		Trees_din <= x"0c004404";
		wait for Clk_period;
		Addr <=  "00010111111101";
		Trees_din <= x"001a180d";
		wait for Clk_period;
		Addr <=  "00010111111110";
		Trees_din <= x"01fa7a04";
		wait for Clk_period;
		Addr <=  "00010111111111";
		Trees_din <= x"ffd1180d";
		wait for Clk_period;
		Addr <=  "00011000000000";
		Trees_din <= x"0006180d";
		wait for Clk_period;
		Addr <=  "00011000000001";
		Trees_din <= x"0028180d";
		wait for Clk_period;
		Addr <=  "00011000000010";
		Trees_din <= x"ffe7180d";
		wait for Clk_period;
		Addr <=  "00011000000011";
		Trees_din <= x"18003004";
		wait for Clk_period;
		Addr <=  "00011000000100";
		Trees_din <= x"001c1829";
		wait for Clk_period;
		Addr <=  "00011000000101";
		Trees_din <= x"04ffce08";
		wait for Clk_period;
		Addr <=  "00011000000110";
		Trees_din <= x"0a018f04";
		wait for Clk_period;
		Addr <=  "00011000000111";
		Trees_din <= x"fff11829";
		wait for Clk_period;
		Addr <=  "00011000001000";
		Trees_din <= x"001f1829";
		wait for Clk_period;
		Addr <=  "00011000001001";
		Trees_din <= x"ffdb1829";
		wait for Clk_period;
		Addr <=  "00011000001010";
		Trees_din <= x"05098d08";
		wait for Clk_period;
		Addr <=  "00011000001011";
		Trees_din <= x"17004504";
		wait for Clk_period;
		Addr <=  "00011000001100";
		Trees_din <= x"ffe1184d";
		wait for Clk_period;
		Addr <=  "00011000001101";
		Trees_din <= x"0009184d";
		wait for Clk_period;
		Addr <=  "00011000001110";
		Trees_din <= x"06fc0e04";
		wait for Clk_period;
		Addr <=  "00011000001111";
		Trees_din <= x"0027184d";
		wait for Clk_period;
		Addr <=  "00011000010000";
		Trees_din <= x"17004104";
		wait for Clk_period;
		Addr <=  "00011000010001";
		Trees_din <= x"0019184d";
		wait for Clk_period;
		Addr <=  "00011000010010";
		Trees_din <= x"ffe7184d";
		wait for Clk_period;
		Addr <=  "00011000010011";
		Trees_din <= x"05085504";
		wait for Clk_period;
		Addr <=  "00011000010100";
		Trees_din <= x"ffec1871";
		wait for Clk_period;
		Addr <=  "00011000010101";
		Trees_din <= x"09fade04";
		wait for Clk_period;
		Addr <=  "00011000010110";
		Trees_din <= x"00201871";
		wait for Clk_period;
		Addr <=  "00011000010111";
		Trees_din <= x"0904f608";
		wait for Clk_period;
		Addr <=  "00011000011000";
		Trees_din <= x"000b0b04";
		wait for Clk_period;
		Addr <=  "00011000011001";
		Trees_din <= x"000a1871";
		wait for Clk_period;
		Addr <=  "00011000011010";
		Trees_din <= x"ffe11871";
		wait for Clk_period;
		Addr <=  "00011000011011";
		Trees_din <= x"00171871";
		wait for Clk_period;
		Addr <=  "00011000011100";
		Trees_din <= x"01027c0c";
		wait for Clk_period;
		Addr <=  "00011000011101";
		Trees_din <= x"10003d04";
		wait for Clk_period;
		Addr <=  "00011000011110";
		Trees_din <= x"ffef188d";
		wait for Clk_period;
		Addr <=  "00011000011111";
		Trees_din <= x"000b0b04";
		wait for Clk_period;
		Addr <=  "00011000100000";
		Trees_din <= x"0029188d";
		wait for Clk_period;
		Addr <=  "00011000100001";
		Trees_din <= x"0001188d";
		wait for Clk_period;
		Addr <=  "00011000100010";
		Trees_din <= x"ffeb188d";
		wait for Clk_period;
		Addr <=  "00011000100011";
		Trees_din <= x"05085504";
		wait for Clk_period;
		Addr <=  "00011000100100";
		Trees_din <= x"ffeb18b1";
		wait for Clk_period;
		Addr <=  "00011000100101";
		Trees_din <= x"03fcf108";
		wait for Clk_period;
		Addr <=  "00011000100110";
		Trees_din <= x"08005304";
		wait for Clk_period;
		Addr <=  "00011000100111";
		Trees_din <= x"000118b1";
		wait for Clk_period;
		Addr <=  "00011000101000";
		Trees_din <= x"002618b1";
		wait for Clk_period;
		Addr <=  "00011000101001";
		Trees_din <= x"18003804";
		wait for Clk_period;
		Addr <=  "00011000101010";
		Trees_din <= x"000e18b1";
		wait for Clk_period;
		Addr <=  "00011000101011";
		Trees_din <= x"ffee18b1";
		wait for Clk_period;
		Addr <=  "00011000101100";
		Trees_din <= x"05098d08";
		wait for Clk_period;
		Addr <=  "00011000101101";
		Trees_din <= x"17004504";
		wait for Clk_period;
		Addr <=  "00011000101110";
		Trees_din <= x"ffe218d5";
		wait for Clk_period;
		Addr <=  "00011000101111";
		Trees_din <= x"000918d5";
		wait for Clk_period;
		Addr <=  "00011000110000";
		Trees_din <= x"06fc0e04";
		wait for Clk_period;
		Addr <=  "00011000110001";
		Trees_din <= x"002318d5";
		wait for Clk_period;
		Addr <=  "00011000110010";
		Trees_din <= x"17004104";
		wait for Clk_period;
		Addr <=  "00011000110011";
		Trees_din <= x"001718d5";
		wait for Clk_period;
		Addr <=  "00011000110100";
		Trees_din <= x"ffeb18d5";
		wait for Clk_period;
		Addr <=  "00011000110101";
		Trees_din <= x"05072404";
		wait for Clk_period;
		Addr <=  "00011000110110";
		Trees_din <= x"ffeb18f9";
		wait for Clk_period;
		Addr <=  "00011000110111";
		Trees_din <= x"03fcf108";
		wait for Clk_period;
		Addr <=  "00011000111000";
		Trees_din <= x"0a013b04";
		wait for Clk_period;
		Addr <=  "00011000111001";
		Trees_din <= x"000018f9";
		wait for Clk_period;
		Addr <=  "00011000111010";
		Trees_din <= x"002618f9";
		wait for Clk_period;
		Addr <=  "00011000111011";
		Trees_din <= x"0a00d404";
		wait for Clk_period;
		Addr <=  "00011000111100";
		Trees_din <= x"000c18f9";
		wait for Clk_period;
		Addr <=  "00011000111101";
		Trees_din <= x"ffed18f9";
		wait for Clk_period;
		Addr <=  "00011000111110";
		Trees_din <= x"18003004";
		wait for Clk_period;
		Addr <=  "00011000111111";
		Trees_din <= x"001a1915";
		wait for Clk_period;
		Addr <=  "00011001000000";
		Trees_din <= x"04ffce08";
		wait for Clk_period;
		Addr <=  "00011001000001";
		Trees_din <= x"0a018f04";
		wait for Clk_period;
		Addr <=  "00011001000010";
		Trees_din <= x"fff31915";
		wait for Clk_period;
		Addr <=  "00011001000011";
		Trees_din <= x"001c1915";
		wait for Clk_period;
		Addr <=  "00011001000100";
		Trees_din <= x"ffde1915";
		wait for Clk_period;
		Addr <=  "00011001000101";
		Trees_din <= x"05098d08";
		wait for Clk_period;
		Addr <=  "00011001000110";
		Trees_din <= x"17004504";
		wait for Clk_period;
		Addr <=  "00011001000111";
		Trees_din <= x"ffe41931";
		wait for Clk_period;
		Addr <=  "00011001001000";
		Trees_din <= x"00071931";
		wait for Clk_period;
		Addr <=  "00011001001001";
		Trees_din <= x"1b01aa04";
		wait for Clk_period;
		Addr <=  "00011001001010";
		Trees_din <= x"001e1931";
		wait for Clk_period;
		Addr <=  "00011001001011";
		Trees_din <= x"fffc1931";
		wait for Clk_period;
		Addr <=  "00011001001100";
		Trees_din <= x"1f040004";
		wait for Clk_period;
		Addr <=  "00011001001101";
		Trees_din <= x"0015194d";
		wait for Clk_period;
		Addr <=  "00011001001110";
		Trees_din <= x"06fc0e04";
		wait for Clk_period;
		Addr <=  "00011001001111";
		Trees_din <= x"001a194d";
		wait for Clk_period;
		Addr <=  "00011001010000";
		Trees_din <= x"0d028004";
		wait for Clk_period;
		Addr <=  "00011001010001";
		Trees_din <= x"ffd8194d";
		wait for Clk_period;
		Addr <=  "00011001010010";
		Trees_din <= x"0004194d";
		wait for Clk_period;
		Addr <=  "00011001010011";
		Trees_din <= x"05085504";
		wait for Clk_period;
		Addr <=  "00011001010100";
		Trees_din <= x"ffed1969";
		wait for Clk_period;
		Addr <=  "00011001010101";
		Trees_din <= x"01f9cc04";
		wait for Clk_period;
		Addr <=  "00011001010110";
		Trees_din <= x"fff71969";
		wait for Clk_period;
		Addr <=  "00011001010111";
		Trees_din <= x"07005604";
		wait for Clk_period;
		Addr <=  "00011001011000";
		Trees_din <= x"00231969";
		wait for Clk_period;
		Addr <=  "00011001011001";
		Trees_din <= x"fffd1969";
		wait for Clk_period;
		Addr <=  "00011001011010";
		Trees_din <= x"0c004504";
		wait for Clk_period;
		Addr <=  "00011001011011";
		Trees_din <= x"00161985";
		wait for Clk_period;
		Addr <=  "00011001011100";
		Trees_din <= x"18003908";
		wait for Clk_period;
		Addr <=  "00011001011101";
		Trees_din <= x"09feb404";
		wait for Clk_period;
		Addr <=  "00011001011110";
		Trees_din <= x"001e1985";
		wait for Clk_period;
		Addr <=  "00011001011111";
		Trees_din <= x"fff31985";
		wait for Clk_period;
		Addr <=  "00011001100000";
		Trees_din <= x"ffe31985";
		wait for Clk_period;
		Addr <=  "00011001100001";
		Trees_din <= x"05098d08";
		wait for Clk_period;
		Addr <=  "00011001100010";
		Trees_din <= x"06fe8904";
		wait for Clk_period;
		Addr <=  "00011001100011";
		Trees_din <= x"ffe619a1";
		wait for Clk_period;
		Addr <=  "00011001100100";
		Trees_din <= x"000219a1";
		wait for Clk_period;
		Addr <=  "00011001100101";
		Trees_din <= x"1b01aa04";
		wait for Clk_period;
		Addr <=  "00011001100110";
		Trees_din <= x"001c19a1";
		wait for Clk_period;
		Addr <=  "00011001100111";
		Trees_din <= x"fffd19a1";
		wait for Clk_period;
		Addr <=  "00011001101000";
		Trees_din <= x"0506f704";
		wait for Clk_period;
		Addr <=  "00011001101001";
		Trees_din <= x"ffeb19c5";
		wait for Clk_period;
		Addr <=  "00011001101010";
		Trees_din <= x"03fcf108";
		wait for Clk_period;
		Addr <=  "00011001101011";
		Trees_din <= x"0a013b04";
		wait for Clk_period;
		Addr <=  "00011001101100";
		Trees_din <= x"fffc19c5";
		wait for Clk_period;
		Addr <=  "00011001101101";
		Trees_din <= x"002519c5";
		wait for Clk_period;
		Addr <=  "00011001101110";
		Trees_din <= x"00087604";
		wait for Clk_period;
		Addr <=  "00011001101111";
		Trees_din <= x"000a19c5";
		wait for Clk_period;
		Addr <=  "00011001110000";
		Trees_din <= x"ffeb19c5";
		wait for Clk_period;
		Addr <=  "00011001110001";
		Trees_din <= x"05098d08";
		wait for Clk_period;
		Addr <=  "00011001110010";
		Trees_din <= x"1b021f04";
		wait for Clk_period;
		Addr <=  "00011001110011";
		Trees_din <= x"ffe819e1";
		wait for Clk_period;
		Addr <=  "00011001110100";
		Trees_din <= x"000319e1";
		wait for Clk_period;
		Addr <=  "00011001110101";
		Trees_din <= x"18003b04";
		wait for Clk_period;
		Addr <=  "00011001110110";
		Trees_din <= x"001a19e1";
		wait for Clk_period;
		Addr <=  "00011001110111";
		Trees_din <= x"fffa19e1";
		wait for Clk_period;
		Addr <=  "00011001111000";
		Trees_din <= x"0a013b08";
		wait for Clk_period;
		Addr <=  "00011001111001";
		Trees_din <= x"0a005a04";
		wait for Clk_period;
		Addr <=  "00011001111010";
		Trees_din <= x"000b19fd";
		wait for Clk_period;
		Addr <=  "00011001111011";
		Trees_din <= x"ffe319fd";
		wait for Clk_period;
		Addr <=  "00011001111100";
		Trees_din <= x"13026d04";
		wait for Clk_period;
		Addr <=  "00011001111101";
		Trees_din <= x"001719fd";
		wait for Clk_period;
		Addr <=  "00011001111110";
		Trees_din <= x"fffc19fd";
		wait for Clk_period;
		Addr <=  "00011001111111";
		Trees_din <= x"05085504";
		wait for Clk_period;
		Addr <=  "00011010000000";
		Trees_din <= x"ffed1a19";
		wait for Clk_period;
		Addr <=  "00011010000001";
		Trees_din <= x"04ffd508";
		wait for Clk_period;
		Addr <=  "00011010000010";
		Trees_din <= x"08005404";
		wait for Clk_period;
		Addr <=  "00011010000011";
		Trees_din <= x"fffc1a19";
		wait for Clk_period;
		Addr <=  "00011010000100";
		Trees_din <= x"00221a19";
		wait for Clk_period;
		Addr <=  "00011010000101";
		Trees_din <= x"fff71a19";
		wait for Clk_period;
		Addr <=  "00011010000110";
		Trees_din <= x"18003004";
		wait for Clk_period;
		Addr <=  "00011010000111";
		Trees_din <= x"00161a35";
		wait for Clk_period;
		Addr <=  "00011010001000";
		Trees_din <= x"04ffce08";
		wait for Clk_period;
		Addr <=  "00011010001001";
		Trees_din <= x"0a018f04";
		wait for Clk_period;
		Addr <=  "00011010001010";
		Trees_din <= x"fff51a35";
		wait for Clk_period;
		Addr <=  "00011010001011";
		Trees_din <= x"00191a35";
		wait for Clk_period;
		Addr <=  "00011010001100";
		Trees_din <= x"ffe01a35";
		wait for Clk_period;
		Addr <=  "00011010001101";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  1
        -----------
		Addr <=  "00000000000000";
		Trees_din <= x"000b0b30";
		wait for Clk_period;
		Addr <=  "00000000000001";
		Trees_din <= x"000a0724";
		wait for Clk_period;
		Addr <=  "00000000000010";
		Trees_din <= x"00087614";
		wait for Clk_period;
		Addr <=  "00000000000011";
		Trees_din <= x"00054904";
		wait for Clk_period;
		Addr <=  "00000000000100";
		Trees_din <= x"ff4d00a5";
		wait for Clk_period;
		Addr <=  "00000000000101";
		Trees_din <= x"03ffbe08";
		wait for Clk_period;
		Addr <=  "00000000000110";
		Trees_din <= x"21000504";
		wait for Clk_period;
		Addr <=  "00000000000111";
		Trees_din <= x"ff5700a5";
		wait for Clk_period;
		Addr <=  "00000000001000";
		Trees_din <= x"ffe500a5";
		wait for Clk_period;
		Addr <=  "00000000001001";
		Trees_din <= x"05012304";
		wait for Clk_period;
		Addr <=  "00000000001010";
		Trees_din <= x"ff9d00a5";
		wait for Clk_period;
		Addr <=  "00000000001011";
		Trees_din <= x"013c00a5";
		wait for Clk_period;
		Addr <=  "00000000001100";
		Trees_din <= x"03fe9a0c";
		wait for Clk_period;
		Addr <=  "00000000001101";
		Trees_din <= x"04001804";
		wait for Clk_period;
		Addr <=  "00000000001110";
		Trees_din <= x"ff5600a5";
		wait for Clk_period;
		Addr <=  "00000000001111";
		Trees_din <= x"03fb9904";
		wait for Clk_period;
		Addr <=  "00000000010000";
		Trees_din <= x"ff9d00a5";
		wait for Clk_period;
		Addr <=  "00000000010001";
		Trees_din <= x"00b200a5";
		wait for Clk_period;
		Addr <=  "00000000010010";
		Trees_din <= x"022400a5";
		wait for Clk_period;
		Addr <=  "00000000010011";
		Trees_din <= x"0507e108";
		wait for Clk_period;
		Addr <=  "00000000010100";
		Trees_din <= x"02083604";
		wait for Clk_period;
		Addr <=  "00000000010101";
		Trees_din <= x"02aa00a5";
		wait for Clk_period;
		Addr <=  "00000000010110";
		Trees_din <= x"ff8100a5";
		wait for Clk_period;
		Addr <=  "00000000010111";
		Trees_din <= x"ff6200a5";
		wait for Clk_period;
		Addr <=  "00000000011000";
		Trees_din <= x"050b070c";
		wait for Clk_period;
		Addr <=  "00000000011001";
		Trees_din <= x"000b6408";
		wait for Clk_period;
		Addr <=  "00000000011010";
		Trees_din <= x"0204f104";
		wait for Clk_period;
		Addr <=  "00000000011011";
		Trees_din <= x"02ca00a5";
		wait for Clk_period;
		Addr <=  "00000000011100";
		Trees_din <= x"000000a5";
		wait for Clk_period;
		Addr <=  "00000000011101";
		Trees_din <= x"042e00a5";
		wait for Clk_period;
		Addr <=  "00000000011110";
		Trees_din <= x"03fcf110";
		wait for Clk_period;
		Addr <=  "00000000011111";
		Trees_din <= x"000c1004";
		wait for Clk_period;
		Addr <=  "00000000100000";
		Trees_din <= x"ff6c00a5";
		wait for Clk_period;
		Addr <=  "00000000100001";
		Trees_din <= x"050d5a08";
		wait for Clk_period;
		Addr <=  "00000000100010";
		Trees_din <= x"04fe6104";
		wait for Clk_period;
		Addr <=  "00000000100011";
		Trees_din <= x"028400a5";
		wait for Clk_period;
		Addr <=  "00000000100100";
		Trees_din <= x"00b200a5";
		wait for Clk_period;
		Addr <=  "00000000100101";
		Trees_din <= x"000000a5";
		wait for Clk_period;
		Addr <=  "00000000100110";
		Trees_din <= x"06fc2004";
		wait for Clk_period;
		Addr <=  "00000000100111";
		Trees_din <= x"00e200a5";
		wait for Clk_period;
		Addr <=  "00000000101000";
		Trees_din <= x"038400a5";
		wait for Clk_period;
		Addr <=  "00000000101001";
		Trees_din <= x"000a072c";
		wait for Clk_period;
		Addr <=  "00000000101010";
		Trees_din <= x"00087618";
		wait for Clk_period;
		Addr <=  "00000000101011";
		Trees_din <= x"00054904";
		wait for Clk_period;
		Addr <=  "00000000101100";
		Trees_din <= x"ff540149";
		wait for Clk_period;
		Addr <=  "00000000101101";
		Trees_din <= x"03ffbe0c";
		wait for Clk_period;
		Addr <=  "00000000101110";
		Trees_din <= x"21000508";
		wait for Clk_period;
		Addr <=  "00000000101111";
		Trees_din <= x"09f74f04";
		wait for Clk_period;
		Addr <=  "00000000110000";
		Trees_din <= x"fff40149";
		wait for Clk_period;
		Addr <=  "00000000110001";
		Trees_din <= x"ff580149";
		wait for Clk_period;
		Addr <=  "00000000110010";
		Trees_din <= x"fff50149";
		wait for Clk_period;
		Addr <=  "00000000110011";
		Trees_din <= x"19009d04";
		wait for Clk_period;
		Addr <=  "00000000110100";
		Trees_din <= x"ff930149";
		wait for Clk_period;
		Addr <=  "00000000110101";
		Trees_din <= x"01370149";
		wait for Clk_period;
		Addr <=  "00000000110110";
		Trees_din <= x"03fe9a0c";
		wait for Clk_period;
		Addr <=  "00000000110111";
		Trees_din <= x"04001804";
		wait for Clk_period;
		Addr <=  "00000000111000";
		Trees_din <= x"ff5e0149";
		wait for Clk_period;
		Addr <=  "00000000111001";
		Trees_din <= x"18003604";
		wait for Clk_period;
		Addr <=  "00000000111010";
		Trees_din <= x"ff9b0149";
		wait for Clk_period;
		Addr <=  "00000000111011";
		Trees_din <= x"00d70149";
		wait for Clk_period;
		Addr <=  "00000000111100";
		Trees_din <= x"02012d04";
		wait for Clk_period;
		Addr <=  "00000000111101";
		Trees_din <= x"01a70149";
		wait for Clk_period;
		Addr <=  "00000000111110";
		Trees_din <= x"002b0149";
		wait for Clk_period;
		Addr <=  "00000000111111";
		Trees_din <= x"000c1024";
		wait for Clk_period;
		Addr <=  "00000001000000";
		Trees_din <= x"050a6c14";
		wait for Clk_period;
		Addr <=  "00000001000001";
		Trees_din <= x"0208360c";
		wait for Clk_period;
		Addr <=  "00000001000010";
		Trees_din <= x"1b002d04";
		wait for Clk_period;
		Addr <=  "00000001000011";
		Trees_din <= x"00450149";
		wait for Clk_period;
		Addr <=  "00000001000100";
		Trees_din <= x"1c002004";
		wait for Clk_period;
		Addr <=  "00000001000101";
		Trees_din <= x"007b0149";
		wait for Clk_period;
		Addr <=  "00000001000110";
		Trees_din <= x"01a20149";
		wait for Clk_period;
		Addr <=  "00000001000111";
		Trees_din <= x"08005904";
		wait for Clk_period;
		Addr <=  "00000001001000";
		Trees_din <= x"ff690149";
		wait for Clk_period;
		Addr <=  "00000001001001";
		Trees_din <= x"002d0149";
		wait for Clk_period;
		Addr <=  "00000001001010";
		Trees_din <= x"03fd0904";
		wait for Clk_period;
		Addr <=  "00000001001011";
		Trees_din <= x"ff630149";
		wait for Clk_period;
		Addr <=  "00000001001100";
		Trees_din <= x"09f96b04";
		wait for Clk_period;
		Addr <=  "00000001001101";
		Trees_din <= x"ff930149";
		wait for Clk_period;
		Addr <=  "00000001001110";
		Trees_din <= x"0b014d04";
		wait for Clk_period;
		Addr <=  "00000001001111";
		Trees_din <= x"00390149";
		wait for Clk_period;
		Addr <=  "00000001010000";
		Trees_din <= x"01800149";
		wait for Clk_period;
		Addr <=  "00000001010001";
		Trees_din <= x"01a80149";
		wait for Clk_period;
		Addr <=  "00000001010010";
		Trees_din <= x"000a0728";
		wait for Clk_period;
		Addr <=  "00000001010011";
		Trees_din <= x"00087618";
		wait for Clk_period;
		Addr <=  "00000001010100";
		Trees_din <= x"00054904";
		wait for Clk_period;
		Addr <=  "00000001010101";
		Trees_din <= x"ff5901fd";
		wait for Clk_period;
		Addr <=  "00000001010110";
		Trees_din <= x"03ffbe0c";
		wait for Clk_period;
		Addr <=  "00000001010111";
		Trees_din <= x"07005c08";
		wait for Clk_period;
		Addr <=  "00000001011000";
		Trees_din <= x"22000104";
		wait for Clk_period;
		Addr <=  "00000001011001";
		Trees_din <= x"ff5d01fd";
		wait for Clk_period;
		Addr <=  "00000001011010";
		Trees_din <= x"000501fd";
		wait for Clk_period;
		Addr <=  "00000001011011";
		Trees_din <= x"000601fd";
		wait for Clk_period;
		Addr <=  "00000001011100";
		Trees_din <= x"00067504";
		wait for Clk_period;
		Addr <=  "00000001011101";
		Trees_din <= x"00f901fd";
		wait for Clk_period;
		Addr <=  "00000001011110";
		Trees_din <= x"ff9501fd";
		wait for Clk_period;
		Addr <=  "00000001011111";
		Trees_din <= x"03fd2804";
		wait for Clk_period;
		Addr <=  "00000001100000";
		Trees_din <= x"ff6401fd";
		wait for Clk_period;
		Addr <=  "00000001100001";
		Trees_din <= x"13028708";
		wait for Clk_period;
		Addr <=  "00000001100010";
		Trees_din <= x"04fe7c04";
		wait for Clk_period;
		Addr <=  "00000001100011";
		Trees_din <= x"002a01fd";
		wait for Clk_period;
		Addr <=  "00000001100100";
		Trees_din <= x"015101fd";
		wait for Clk_period;
		Addr <=  "00000001100101";
		Trees_din <= x"ff9201fd";
		wait for Clk_period;
		Addr <=  "00000001100110";
		Trees_din <= x"050d5a24";
		wait for Clk_period;
		Addr <=  "00000001100111";
		Trees_din <= x"000bb818";
		wait for Clk_period;
		Addr <=  "00000001101000";
		Trees_din <= x"03fdbf10";
		wait for Clk_period;
		Addr <=  "00000001101001";
		Trees_din <= x"01fd8208";
		wait for Clk_period;
		Addr <=  "00000001101010";
		Trees_din <= x"1c003104";
		wait for Clk_period;
		Addr <=  "00000001101011";
		Trees_din <= x"00c301fd";
		wait for Clk_period;
		Addr <=  "00000001101100";
		Trees_din <= x"ff9601fd";
		wait for Clk_period;
		Addr <=  "00000001101101";
		Trees_din <= x"020d6204";
		wait for Clk_period;
		Addr <=  "00000001101110";
		Trees_din <= x"00f701fd";
		wait for Clk_period;
		Addr <=  "00000001101111";
		Trees_din <= x"ff9801fd";
		wait for Clk_period;
		Addr <=  "00000001110000";
		Trees_din <= x"0f02af04";
		wait for Clk_period;
		Addr <=  "00000001110001";
		Trees_din <= x"014c01fd";
		wait for Clk_period;
		Addr <=  "00000001110010";
		Trees_din <= x"000001fd";
		wait for Clk_period;
		Addr <=  "00000001110011";
		Trees_din <= x"03f9ea04";
		wait for Clk_period;
		Addr <=  "00000001110100";
		Trees_din <= x"005101fd";
		wait for Clk_period;
		Addr <=  "00000001110101";
		Trees_din <= x"04078904";
		wait for Clk_period;
		Addr <=  "00000001110110";
		Trees_din <= x"013101fd";
		wait for Clk_period;
		Addr <=  "00000001110111";
		Trees_din <= x"007d01fd";
		wait for Clk_period;
		Addr <=  "00000001111000";
		Trees_din <= x"03fd0908";
		wait for Clk_period;
		Addr <=  "00000001111001";
		Trees_din <= x"1403c604";
		wait for Clk_period;
		Addr <=  "00000001111010";
		Trees_din <= x"ff6901fd";
		wait for Clk_period;
		Addr <=  "00000001111011";
		Trees_din <= x"003d01fd";
		wait for Clk_period;
		Addr <=  "00000001111100";
		Trees_din <= x"0f028704";
		wait for Clk_period;
		Addr <=  "00000001111101";
		Trees_din <= x"011201fd";
		wait for Clk_period;
		Addr <=  "00000001111110";
		Trees_din <= x"000401fd";
		wait for Clk_period;
		Addr <=  "00000001111111";
		Trees_din <= x"000a0728";
		wait for Clk_period;
		Addr <=  "00000010000000";
		Trees_din <= x"0007ff14";
		wait for Clk_period;
		Addr <=  "00000010000001";
		Trees_din <= x"00054904";
		wait for Clk_period;
		Addr <=  "00000010000010";
		Trees_din <= x"ff5c02a9";
		wait for Clk_period;
		Addr <=  "00000010000011";
		Trees_din <= x"03ffbe08";
		wait for Clk_period;
		Addr <=  "00000010000100";
		Trees_din <= x"21000504";
		wait for Clk_period;
		Addr <=  "00000010000101";
		Trees_din <= x"ff6202a9";
		wait for Clk_period;
		Addr <=  "00000010000110";
		Trees_din <= x"003002a9";
		wait for Clk_period;
		Addr <=  "00000010000111";
		Trees_din <= x"00067504";
		wait for Clk_period;
		Addr <=  "00000010001000";
		Trees_din <= x"00c602a9";
		wait for Clk_period;
		Addr <=  "00000010001001";
		Trees_din <= x"ff9b02a9";
		wait for Clk_period;
		Addr <=  "00000010001010";
		Trees_din <= x"03fd2804";
		wait for Clk_period;
		Addr <=  "00000010001011";
		Trees_din <= x"ff6602a9";
		wait for Clk_period;
		Addr <=  "00000010001100";
		Trees_din <= x"04fecb08";
		wait for Clk_period;
		Addr <=  "00000010001101";
		Trees_din <= x"1b030204";
		wait for Clk_period;
		Addr <=  "00000010001110";
		Trees_din <= x"ff8c02a9";
		wait for Clk_period;
		Addr <=  "00000010001111";
		Trees_din <= x"002b02a9";
		wait for Clk_period;
		Addr <=  "00000010010000";
		Trees_din <= x"05fb6c04";
		wait for Clk_period;
		Addr <=  "00000010010001";
		Trees_din <= x"002f02a9";
		wait for Clk_period;
		Addr <=  "00000010010010";
		Trees_din <= x"013002a9";
		wait for Clk_period;
		Addr <=  "00000010010011";
		Trees_din <= x"000c1024";
		wait for Clk_period;
		Addr <=  "00000010010100";
		Trees_din <= x"03fdbf18";
		wait for Clk_period;
		Addr <=  "00000010010101";
		Trees_din <= x"050a6c10";
		wait for Clk_period;
		Addr <=  "00000010010110";
		Trees_din <= x"0206da08";
		wait for Clk_period;
		Addr <=  "00000010010111";
		Trees_din <= x"1b002d04";
		wait for Clk_period;
		Addr <=  "00000010011000";
		Trees_din <= x"ff8a02a9";
		wait for Clk_period;
		Addr <=  "00000010011001";
		Trees_din <= x"00c502a9";
		wait for Clk_period;
		Addr <=  "00000010011010";
		Trees_din <= x"04013a04";
		wait for Clk_period;
		Addr <=  "00000010011011";
		Trees_din <= x"ff6e02a9";
		wait for Clk_period;
		Addr <=  "00000010011100";
		Trees_din <= x"003902a9";
		wait for Clk_period;
		Addr <=  "00000010011101";
		Trees_din <= x"1505d604";
		wait for Clk_period;
		Addr <=  "00000010011110";
		Trees_din <= x"ff6a02a9";
		wait for Clk_period;
		Addr <=  "00000010011111";
		Trees_din <= x"00a902a9";
		wait for Clk_period;
		Addr <=  "00000010100000";
		Trees_din <= x"1603f208";
		wait for Clk_period;
		Addr <=  "00000010100001";
		Trees_din <= x"0b043e04";
		wait for Clk_period;
		Addr <=  "00000010100010";
		Trees_din <= x"010a02a9";
		wait for Clk_period;
		Addr <=  "00000010100011";
		Trees_din <= x"002802a9";
		wait for Clk_period;
		Addr <=  "00000010100100";
		Trees_din <= x"000002a9";
		wait for Clk_period;
		Addr <=  "00000010100101";
		Trees_din <= x"03f9ea04";
		wait for Clk_period;
		Addr <=  "00000010100110";
		Trees_din <= x"002602a9";
		wait for Clk_period;
		Addr <=  "00000010100111";
		Trees_din <= x"04078904";
		wait for Clk_period;
		Addr <=  "00000010101000";
		Trees_din <= x"00f802a9";
		wait for Clk_period;
		Addr <=  "00000010101001";
		Trees_din <= x"006702a9";
		wait for Clk_period;
		Addr <=  "00000010101010";
		Trees_din <= x"000a0728";
		wait for Clk_period;
		Addr <=  "00000010101011";
		Trees_din <= x"0007ff14";
		wait for Clk_period;
		Addr <=  "00000010101100";
		Trees_din <= x"00054904";
		wait for Clk_period;
		Addr <=  "00000010101101";
		Trees_din <= x"ff5f0385";
		wait for Clk_period;
		Addr <=  "00000010101110";
		Trees_din <= x"03ffbe08";
		wait for Clk_period;
		Addr <=  "00000010101111";
		Trees_din <= x"21000504";
		wait for Clk_period;
		Addr <=  "00000010110000";
		Trees_din <= x"ff660385";
		wait for Clk_period;
		Addr <=  "00000010110001";
		Trees_din <= x"00320385";
		wait for Clk_period;
		Addr <=  "00000010110010";
		Trees_din <= x"19009d04";
		wait for Clk_period;
		Addr <=  "00000010110011";
		Trees_din <= x"ff9f0385";
		wait for Clk_period;
		Addr <=  "00000010110100";
		Trees_din <= x"00a80385";
		wait for Clk_period;
		Addr <=  "00000010110101";
		Trees_din <= x"03fd2804";
		wait for Clk_period;
		Addr <=  "00000010110110";
		Trees_din <= x"ff6b0385";
		wait for Clk_period;
		Addr <=  "00000010110111";
		Trees_din <= x"04fecb08";
		wait for Clk_period;
		Addr <=  "00000010111000";
		Trees_din <= x"1b030204";
		wait for Clk_period;
		Addr <=  "00000010111001";
		Trees_din <= x"ff930385";
		wait for Clk_period;
		Addr <=  "00000010111010";
		Trees_din <= x"00270385";
		wait for Clk_period;
		Addr <=  "00000010111011";
		Trees_din <= x"18003604";
		wait for Clk_period;
		Addr <=  "00000010111100";
		Trees_din <= x"00340385";
		wait for Clk_period;
		Addr <=  "00000010111101";
		Trees_din <= x"010c0385";
		wait for Clk_period;
		Addr <=  "00000010111110";
		Trees_din <= x"000c102c";
		wait for Clk_period;
		Addr <=  "00000010111111";
		Trees_din <= x"03fdbf20";
		wait for Clk_period;
		Addr <=  "00000011000000";
		Trees_din <= x"05072410";
		wait for Clk_period;
		Addr <=  "00000011000001";
		Trees_din <= x"0206da08";
		wait for Clk_period;
		Addr <=  "00000011000010";
		Trees_din <= x"04007104";
		wait for Clk_period;
		Addr <=  "00000011000011";
		Trees_din <= x"00c80385";
		wait for Clk_period;
		Addr <=  "00000011000100";
		Trees_din <= x"ffb70385";
		wait for Clk_period;
		Addr <=  "00000011000101";
		Trees_din <= x"04013a04";
		wait for Clk_period;
		Addr <=  "00000011000110";
		Trees_din <= x"ff7a0385";
		wait for Clk_period;
		Addr <=  "00000011000111";
		Trees_din <= x"003d0385";
		wait for Clk_period;
		Addr <=  "00000011001000";
		Trees_din <= x"13fb2408";
		wait for Clk_period;
		Addr <=  "00000011001001";
		Trees_din <= x"0c00af04";
		wait for Clk_period;
		Addr <=  "00000011001010";
		Trees_din <= x"ffa70385";
		wait for Clk_period;
		Addr <=  "00000011001011";
		Trees_din <= x"00b10385";
		wait for Clk_period;
		Addr <=  "00000011001100";
		Trees_din <= x"08004504";
		wait for Clk_period;
		Addr <=  "00000011001101";
		Trees_din <= x"005b0385";
		wait for Clk_period;
		Addr <=  "00000011001110";
		Trees_din <= x"ff540385";
		wait for Clk_period;
		Addr <=  "00000011001111";
		Trees_din <= x"1603f208";
		wait for Clk_period;
		Addr <=  "00000011010000";
		Trees_din <= x"0b043e04";
		wait for Clk_period;
		Addr <=  "00000011010001";
		Trees_din <= x"00e00385";
		wait for Clk_period;
		Addr <=  "00000011010010";
		Trees_din <= x"00170385";
		wait for Clk_period;
		Addr <=  "00000011010011";
		Trees_din <= x"fff80385";
		wait for Clk_period;
		Addr <=  "00000011010100";
		Trees_din <= x"050d5a10";
		wait for Clk_period;
		Addr <=  "00000011010101";
		Trees_din <= x"03f9ea04";
		wait for Clk_period;
		Addr <=  "00000011010110";
		Trees_din <= x"00340385";
		wait for Clk_period;
		Addr <=  "00000011010111";
		Trees_din <= x"04078908";
		wait for Clk_period;
		Addr <=  "00000011011000";
		Trees_din <= x"05085504";
		wait for Clk_period;
		Addr <=  "00000011011001";
		Trees_din <= x"00d90385";
		wait for Clk_period;
		Addr <=  "00000011011010";
		Trees_din <= x"00bd0385";
		wait for Clk_period;
		Addr <=  "00000011011011";
		Trees_din <= x"00510385";
		wait for Clk_period;
		Addr <=  "00000011011100";
		Trees_din <= x"13fadb04";
		wait for Clk_period;
		Addr <=  "00000011011101";
		Trees_din <= x"ff7f0385";
		wait for Clk_period;
		Addr <=  "00000011011110";
		Trees_din <= x"15028704";
		wait for Clk_period;
		Addr <=  "00000011011111";
		Trees_din <= x"00da0385";
		wait for Clk_period;
		Addr <=  "00000011100000";
		Trees_din <= x"00110385";
		wait for Clk_period;
		Addr <=  "00000011100001";
		Trees_din <= x"000a0728";
		wait for Clk_period;
		Addr <=  "00000011100010";
		Trees_din <= x"0007ff14";
		wait for Clk_period;
		Addr <=  "00000011100011";
		Trees_din <= x"00054904";
		wait for Clk_period;
		Addr <=  "00000011100100";
		Trees_din <= x"ff610471";
		wait for Clk_period;
		Addr <=  "00000011100101";
		Trees_din <= x"03ffbe08";
		wait for Clk_period;
		Addr <=  "00000011100110";
		Trees_din <= x"22000104";
		wait for Clk_period;
		Addr <=  "00000011100111";
		Trees_din <= x"ff6a0471";
		wait for Clk_period;
		Addr <=  "00000011101000";
		Trees_din <= x"003c0471";
		wait for Clk_period;
		Addr <=  "00000011101001";
		Trees_din <= x"19009d04";
		wait for Clk_period;
		Addr <=  "00000011101010";
		Trees_din <= x"ffa50471";
		wait for Clk_period;
		Addr <=  "00000011101011";
		Trees_din <= x"008d0471";
		wait for Clk_period;
		Addr <=  "00000011101100";
		Trees_din <= x"03fd2804";
		wait for Clk_period;
		Addr <=  "00000011101101";
		Trees_din <= x"ff700471";
		wait for Clk_period;
		Addr <=  "00000011101110";
		Trees_din <= x"04fecb08";
		wait for Clk_period;
		Addr <=  "00000011101111";
		Trees_din <= x"1000e704";
		wait for Clk_period;
		Addr <=  "00000011110000";
		Trees_din <= x"00210471";
		wait for Clk_period;
		Addr <=  "00000011110001";
		Trees_din <= x"ff9a0471";
		wait for Clk_period;
		Addr <=  "00000011110010";
		Trees_din <= x"18003604";
		wait for Clk_period;
		Addr <=  "00000011110011";
		Trees_din <= x"00290471";
		wait for Clk_period;
		Addr <=  "00000011110100";
		Trees_din <= x"00e20471";
		wait for Clk_period;
		Addr <=  "00000011110101";
		Trees_din <= x"000c1028";
		wait for Clk_period;
		Addr <=  "00000011110110";
		Trees_din <= x"03fdbf18";
		wait for Clk_period;
		Addr <=  "00000011110111";
		Trees_din <= x"1e007810";
		wait for Clk_period;
		Addr <=  "00000011111000";
		Trees_din <= x"02ffab08";
		wait for Clk_period;
		Addr <=  "00000011111001";
		Trees_din <= x"14030604";
		wait for Clk_period;
		Addr <=  "00000011111010";
		Trees_din <= x"ff4c0471";
		wait for Clk_period;
		Addr <=  "00000011111011";
		Trees_din <= x"004c0471";
		wait for Clk_period;
		Addr <=  "00000011111100";
		Trees_din <= x"09043d04";
		wait for Clk_period;
		Addr <=  "00000011111101";
		Trees_din <= x"00ae0471";
		wait for Clk_period;
		Addr <=  "00000011111110";
		Trees_din <= x"ffcc0471";
		wait for Clk_period;
		Addr <=  "00000011111111";
		Trees_din <= x"0e014804";
		wait for Clk_period;
		Addr <=  "00000100000000";
		Trees_din <= x"ff6a0471";
		wait for Clk_period;
		Addr <=  "00000100000001";
		Trees_din <= x"003f0471";
		wait for Clk_period;
		Addr <=  "00000100000010";
		Trees_din <= x"09faf108";
		wait for Clk_period;
		Addr <=  "00000100000011";
		Trees_din <= x"03fe8c04";
		wait for Clk_period;
		Addr <=  "00000100000100";
		Trees_din <= x"00890471";
		wait for Clk_period;
		Addr <=  "00000100000101";
		Trees_din <= x"ffc20471";
		wait for Clk_period;
		Addr <=  "00000100000110";
		Trees_din <= x"0905c704";
		wait for Clk_period;
		Addr <=  "00000100000111";
		Trees_din <= x"00ce0471";
		wait for Clk_period;
		Addr <=  "00000100001000";
		Trees_din <= x"00380471";
		wait for Clk_period;
		Addr <=  "00000100001001";
		Trees_din <= x"05085508";
		wait for Clk_period;
		Addr <=  "00000100001010";
		Trees_din <= x"04078904";
		wait for Clk_period;
		Addr <=  "00000100001011";
		Trees_din <= x"00c50471";
		wait for Clk_period;
		Addr <=  "00000100001100";
		Trees_din <= x"00410471";
		wait for Clk_period;
		Addr <=  "00000100001101";
		Trees_din <= x"08005810";
		wait for Clk_period;
		Addr <=  "00000100001110";
		Trees_din <= x"09f76208";
		wait for Clk_period;
		Addr <=  "00000100001111";
		Trees_din <= x"0a015404";
		wait for Clk_period;
		Addr <=  "00000100010000";
		Trees_din <= x"00720471";
		wait for Clk_period;
		Addr <=  "00000100010001";
		Trees_din <= x"ff7e0471";
		wait for Clk_period;
		Addr <=  "00000100010010";
		Trees_din <= x"1200b304";
		wait for Clk_period;
		Addr <=  "00000100010011";
		Trees_din <= x"00c40471";
		wait for Clk_period;
		Addr <=  "00000100010100";
		Trees_din <= x"002d0471";
		wait for Clk_period;
		Addr <=  "00000100010101";
		Trees_din <= x"03fc8808";
		wait for Clk_period;
		Addr <=  "00000100010110";
		Trees_din <= x"14031b04";
		wait for Clk_period;
		Addr <=  "00000100010111";
		Trees_din <= x"ff1d0471";
		wait for Clk_period;
		Addr <=  "00000100011000";
		Trees_din <= x"000c0471";
		wait for Clk_period;
		Addr <=  "00000100011001";
		Trees_din <= x"11036f04";
		wait for Clk_period;
		Addr <=  "00000100011010";
		Trees_din <= x"00a80471";
		wait for Clk_period;
		Addr <=  "00000100011011";
		Trees_din <= x"000e0471";
		wait for Clk_period;
		Addr <=  "00000100011100";
		Trees_din <= x"000b0b38";
		wait for Clk_period;
		Addr <=  "00000100011101";
		Trees_din <= x"0007ff14";
		wait for Clk_period;
		Addr <=  "00000100011110";
		Trees_din <= x"00054904";
		wait for Clk_period;
		Addr <=  "00000100011111";
		Trees_din <= x"ff63055d";
		wait for Clk_period;
		Addr <=  "00000100100000";
		Trees_din <= x"11035308";
		wait for Clk_period;
		Addr <=  "00000100100001";
		Trees_din <= x"1b036404";
		wait for Clk_period;
		Addr <=  "00000100100010";
		Trees_din <= x"ff6d055d";
		wait for Clk_period;
		Addr <=  "00000100100011";
		Trees_din <= x"0001055d";
		wait for Clk_period;
		Addr <=  "00000100100100";
		Trees_din <= x"1b020004";
		wait for Clk_period;
		Addr <=  "00000100100101";
		Trees_din <= x"0096055d";
		wait for Clk_period;
		Addr <=  "00000100100110";
		Trees_din <= x"ffa1055d";
		wait for Clk_period;
		Addr <=  "00000100100111";
		Trees_din <= x"03ff4c1c";
		wait for Clk_period;
		Addr <=  "00000100101000";
		Trees_din <= x"15048210";
		wait for Clk_period;
		Addr <=  "00000100101001";
		Trees_din <= x"08005608";
		wait for Clk_period;
		Addr <=  "00000100101010";
		Trees_din <= x"0c028704";
		wait for Clk_period;
		Addr <=  "00000100101011";
		Trees_din <= x"ff55055d";
		wait for Clk_period;
		Addr <=  "00000100101100";
		Trees_din <= x"fff9055d";
		wait for Clk_period;
		Addr <=  "00000100101101";
		Trees_din <= x"0507e104";
		wait for Clk_period;
		Addr <=  "00000100101110";
		Trees_din <= x"0054055d";
		wait for Clk_period;
		Addr <=  "00000100101111";
		Trees_din <= x"ff8d055d";
		wait for Clk_period;
		Addr <=  "00000100110000";
		Trees_din <= x"03fcbe04";
		wait for Clk_period;
		Addr <=  "00000100110001";
		Trees_din <= x"ff9d055d";
		wait for Clk_period;
		Addr <=  "00000100110010";
		Trees_din <= x"08005204";
		wait for Clk_period;
		Addr <=  "00000100110011";
		Trees_din <= x"00c8055d";
		wait for Clk_period;
		Addr <=  "00000100110100";
		Trees_din <= x"002d055d";
		wait for Clk_period;
		Addr <=  "00000100110101";
		Trees_din <= x"1f040004";
		wait for Clk_period;
		Addr <=  "00000100110110";
		Trees_din <= x"000f055d";
		wait for Clk_period;
		Addr <=  "00000100110111";
		Trees_din <= x"00b9055d";
		wait for Clk_period;
		Addr <=  "00000100111000";
		Trees_din <= x"05085514";
		wait for Clk_period;
		Addr <=  "00000100111001";
		Trees_din <= x"04078910";
		wait for Clk_period;
		Addr <=  "00000100111010";
		Trees_din <= x"000c100c";
		wait for Clk_period;
		Addr <=  "00000100111011";
		Trees_din <= x"0ef86f04";
		wait for Clk_period;
		Addr <=  "00000100111100";
		Trees_din <= x"ffb3055d";
		wait for Clk_period;
		Addr <=  "00000100111101";
		Trees_din <= x"0206da04";
		wait for Clk_period;
		Addr <=  "00000100111110";
		Trees_din <= x"00ac055d";
		wait for Clk_period;
		Addr <=  "00000100111111";
		Trees_din <= x"fffb055d";
		wait for Clk_period;
		Addr <=  "00000101000000";
		Trees_din <= x"00b8055d";
		wait for Clk_period;
		Addr <=  "00000101000001";
		Trees_din <= x"0034055d";
		wait for Clk_period;
		Addr <=  "00000101000010";
		Trees_din <= x"0800581c";
		wait for Clk_period;
		Addr <=  "00000101000011";
		Trees_din <= x"09f96b10";
		wait for Clk_period;
		Addr <=  "00000101000100";
		Trees_din <= x"12009608";
		wait for Clk_period;
		Addr <=  "00000101000101";
		Trees_din <= x"0a015404";
		wait for Clk_period;
		Addr <=  "00000101000110";
		Trees_din <= x"0021055d";
		wait for Clk_period;
		Addr <=  "00000101000111";
		Trees_din <= x"ff52055d";
		wait for Clk_period;
		Addr <=  "00000101001000";
		Trees_din <= x"06fc9204";
		wait for Clk_period;
		Addr <=  "00000101001001";
		Trees_din <= x"001d055d";
		wait for Clk_period;
		Addr <=  "00000101001010";
		Trees_din <= x"008c055d";
		wait for Clk_period;
		Addr <=  "00000101001011";
		Trees_din <= x"03fcf108";
		wait for Clk_period;
		Addr <=  "00000101001100";
		Trees_din <= x"000c1004";
		wait for Clk_period;
		Addr <=  "00000101001101";
		Trees_din <= x"ffb7055d";
		wait for Clk_period;
		Addr <=  "00000101001110";
		Trees_din <= x"0095055d";
		wait for Clk_period;
		Addr <=  "00000101001111";
		Trees_din <= x"00c0055d";
		wait for Clk_period;
		Addr <=  "00000101010000";
		Trees_din <= x"03fc8808";
		wait for Clk_period;
		Addr <=  "00000101010001";
		Trees_din <= x"14031b04";
		wait for Clk_period;
		Addr <=  "00000101010010";
		Trees_din <= x"ff3f055d";
		wait for Clk_period;
		Addr <=  "00000101010011";
		Trees_din <= x"0008055d";
		wait for Clk_period;
		Addr <=  "00000101010100";
		Trees_din <= x"11036f04";
		wait for Clk_period;
		Addr <=  "00000101010101";
		Trees_din <= x"0098055d";
		wait for Clk_period;
		Addr <=  "00000101010110";
		Trees_din <= x"0006055d";
		wait for Clk_period;
		Addr <=  "00000101010111";
		Trees_din <= x"000b0b38";
		wait for Clk_period;
		Addr <=  "00000101011000";
		Trees_din <= x"0007ff14";
		wait for Clk_period;
		Addr <=  "00000101011001";
		Trees_din <= x"00054904";
		wait for Clk_period;
		Addr <=  "00000101011010";
		Trees_din <= x"ff640639";
		wait for Clk_period;
		Addr <=  "00000101011011";
		Trees_din <= x"11035308";
		wait for Clk_period;
		Addr <=  "00000101011100";
		Trees_din <= x"1b036404";
		wait for Clk_period;
		Addr <=  "00000101011101";
		Trees_din <= x"ff720639";
		wait for Clk_period;
		Addr <=  "00000101011110";
		Trees_din <= x"00030639";
		wait for Clk_period;
		Addr <=  "00000101011111";
		Trees_din <= x"18003704";
		wait for Clk_period;
		Addr <=  "00000101100000";
		Trees_din <= x"008a0639";
		wait for Clk_period;
		Addr <=  "00000101100001";
		Trees_din <= x"ffa80639";
		wait for Clk_period;
		Addr <=  "00000101100010";
		Trees_din <= x"03ff4c1c";
		wait for Clk_period;
		Addr <=  "00000101100011";
		Trees_din <= x"15048210";
		wait for Clk_period;
		Addr <=  "00000101100100";
		Trees_din <= x"08005608";
		wait for Clk_period;
		Addr <=  "00000101100101";
		Trees_din <= x"0c028704";
		wait for Clk_period;
		Addr <=  "00000101100110";
		Trees_din <= x"ff570639";
		wait for Clk_period;
		Addr <=  "00000101100111";
		Trees_din <= x"fffb0639";
		wait for Clk_period;
		Addr <=  "00000101101000";
		Trees_din <= x"0507e104";
		wait for Clk_period;
		Addr <=  "00000101101001";
		Trees_din <= x"00450639";
		wait for Clk_period;
		Addr <=  "00000101101010";
		Trees_din <= x"ff950639";
		wait for Clk_period;
		Addr <=  "00000101101011";
		Trees_din <= x"03fcbe04";
		wait for Clk_period;
		Addr <=  "00000101101100";
		Trees_din <= x"ffa40639";
		wait for Clk_period;
		Addr <=  "00000101101101";
		Trees_din <= x"08005204";
		wait for Clk_period;
		Addr <=  "00000101101110";
		Trees_din <= x"00ac0639";
		wait for Clk_period;
		Addr <=  "00000101101111";
		Trees_din <= x"00260639";
		wait for Clk_period;
		Addr <=  "00000101110000";
		Trees_din <= x"1f040004";
		wait for Clk_period;
		Addr <=  "00000101110001";
		Trees_din <= x"00030639";
		wait for Clk_period;
		Addr <=  "00000101110010";
		Trees_din <= x"00a60639";
		wait for Clk_period;
		Addr <=  "00000101110011";
		Trees_din <= x"000e0628";
		wait for Clk_period;
		Addr <=  "00000101110100";
		Trees_din <= x"03fd4618";
		wait for Clk_period;
		Addr <=  "00000101110101";
		Trees_din <= x"01fd3510";
		wait for Clk_period;
		Addr <=  "00000101110110";
		Trees_din <= x"12009608";
		wait for Clk_period;
		Addr <=  "00000101110111";
		Trees_din <= x"1e006b04";
		wait for Clk_period;
		Addr <=  "00000101111000";
		Trees_din <= x"ff380639";
		wait for Clk_period;
		Addr <=  "00000101111001";
		Trees_din <= x"00290639";
		wait for Clk_period;
		Addr <=  "00000101111010";
		Trees_din <= x"050c4e04";
		wait for Clk_period;
		Addr <=  "00000101111011";
		Trees_din <= x"00980639";
		wait for Clk_period;
		Addr <=  "00000101111100";
		Trees_din <= x"ffb10639";
		wait for Clk_period;
		Addr <=  "00000101111101";
		Trees_din <= x"09055904";
		wait for Clk_period;
		Addr <=  "00000101111110";
		Trees_din <= x"00a80639";
		wait for Clk_period;
		Addr <=  "00000101111111";
		Trees_din <= x"ffed0639";
		wait for Clk_period;
		Addr <=  "00000110000000";
		Trees_din <= x"0d001104";
		wait for Clk_period;
		Addr <=  "00000110000001";
		Trees_din <= x"fffd0639";
		wait for Clk_period;
		Addr <=  "00000110000010";
		Trees_din <= x"02faa208";
		wait for Clk_period;
		Addr <=  "00000110000011";
		Trees_din <= x"0f02a904";
		wait for Clk_period;
		Addr <=  "00000110000100";
		Trees_din <= x"00990639";
		wait for Clk_period;
		Addr <=  "00000110000101";
		Trees_din <= x"ff8d0639";
		wait for Clk_period;
		Addr <=  "00000110000110";
		Trees_din <= x"00af0639";
		wait for Clk_period;
		Addr <=  "00000110000111";
		Trees_din <= x"0407890c";
		wait for Clk_period;
		Addr <=  "00000110001000";
		Trees_din <= x"03fafa08";
		wait for Clk_period;
		Addr <=  "00000110001001";
		Trees_din <= x"04fe2204";
		wait for Clk_period;
		Addr <=  "00000110001010";
		Trees_din <= x"ffe90639";
		wait for Clk_period;
		Addr <=  "00000110001011";
		Trees_din <= x"00810639";
		wait for Clk_period;
		Addr <=  "00000110001100";
		Trees_din <= x"00af0639";
		wait for Clk_period;
		Addr <=  "00000110001101";
		Trees_din <= x"002c0639";
		wait for Clk_period;
		Addr <=  "00000110001110";
		Trees_din <= x"000b0b2c";
		wait for Clk_period;
		Addr <=  "00000110001111";
		Trees_din <= x"00054904";
		wait for Clk_period;
		Addr <=  "00000110010000";
		Trees_din <= x"ff650715";
		wait for Clk_period;
		Addr <=  "00000110010001";
		Trees_din <= x"03ff4c18";
		wait for Clk_period;
		Addr <=  "00000110010010";
		Trees_din <= x"04fee808";
		wait for Clk_period;
		Addr <=  "00000110010011";
		Trees_din <= x"000a8004";
		wait for Clk_period;
		Addr <=  "00000110010100";
		Trees_din <= x"ff700715";
		wait for Clk_period;
		Addr <=  "00000110010101";
		Trees_din <= x"ffef0715";
		wait for Clk_period;
		Addr <=  "00000110010110";
		Trees_din <= x"15048208";
		wait for Clk_period;
		Addr <=  "00000110010111";
		Trees_din <= x"08005404";
		wait for Clk_period;
		Addr <=  "00000110011000";
		Trees_din <= x"ff710715";
		wait for Clk_period;
		Addr <=  "00000110011001";
		Trees_din <= x"00000715";
		wait for Clk_period;
		Addr <=  "00000110011010";
		Trees_din <= x"01fc4704";
		wait for Clk_period;
		Addr <=  "00000110011011";
		Trees_din <= x"00c30715";
		wait for Clk_period;
		Addr <=  "00000110011100";
		Trees_din <= x"fffd0715";
		wait for Clk_period;
		Addr <=  "00000110011101";
		Trees_din <= x"1f040004";
		wait for Clk_period;
		Addr <=  "00000110011110";
		Trees_din <= x"ffce0715";
		wait for Clk_period;
		Addr <=  "00000110011111";
		Trees_din <= x"0007ff08";
		wait for Clk_period;
		Addr <=  "00000110100000";
		Trees_din <= x"01fa1804";
		wait for Clk_period;
		Addr <=  "00000110100001";
		Trees_din <= x"004c0715";
		wait for Clk_period;
		Addr <=  "00000110100010";
		Trees_din <= x"fff20715";
		wait for Clk_period;
		Addr <=  "00000110100011";
		Trees_din <= x"00990715";
		wait for Clk_period;
		Addr <=  "00000110100100";
		Trees_din <= x"000e062c";
		wait for Clk_period;
		Addr <=  "00000110100101";
		Trees_din <= x"03fd461c";
		wait for Clk_period;
		Addr <=  "00000110100110";
		Trees_din <= x"0904f30c";
		wait for Clk_period;
		Addr <=  "00000110100111";
		Trees_din <= x"03fd3608";
		wait for Clk_period;
		Addr <=  "00000110101000";
		Trees_din <= x"02feff04";
		wait for Clk_period;
		Addr <=  "00000110101001";
		Trees_din <= x"ffe00715";
		wait for Clk_period;
		Addr <=  "00000110101010";
		Trees_din <= x"00900715";
		wait for Clk_period;
		Addr <=  "00000110101011";
		Trees_din <= x"ff7f0715";
		wait for Clk_period;
		Addr <=  "00000110101100";
		Trees_din <= x"05072408";
		wait for Clk_period;
		Addr <=  "00000110101101";
		Trees_din <= x"14036304";
		wait for Clk_period;
		Addr <=  "00000110101110";
		Trees_din <= x"00770715";
		wait for Clk_period;
		Addr <=  "00000110101111";
		Trees_din <= x"fff90715";
		wait for Clk_period;
		Addr <=  "00000110110000";
		Trees_din <= x"0c00da04";
		wait for Clk_period;
		Addr <=  "00000110110001";
		Trees_din <= x"ff4b0715";
		wait for Clk_period;
		Addr <=  "00000110110010";
		Trees_din <= x"ffdc0715";
		wait for Clk_period;
		Addr <=  "00000110110011";
		Trees_din <= x"1403fe0c";
		wait for Clk_period;
		Addr <=  "00000110110100";
		Trees_din <= x"02faa208";
		wait for Clk_period;
		Addr <=  "00000110110101";
		Trees_din <= x"1b01b104";
		wait for Clk_period;
		Addr <=  "00000110110110";
		Trees_din <= x"00990715";
		wait for Clk_period;
		Addr <=  "00000110110111";
		Trees_din <= x"ff9b0715";
		wait for Clk_period;
		Addr <=  "00000110111000";
		Trees_din <= x"00a70715";
		wait for Clk_period;
		Addr <=  "00000110111001";
		Trees_din <= x"fff50715";
		wait for Clk_period;
		Addr <=  "00000110111010";
		Trees_din <= x"04078914";
		wait for Clk_period;
		Addr <=  "00000110111011";
		Trees_din <= x"0508d704";
		wait for Clk_period;
		Addr <=  "00000110111100";
		Trees_din <= x"00a90715";
		wait for Clk_period;
		Addr <=  "00000110111101";
		Trees_din <= x"1d009308";
		wait for Clk_period;
		Addr <=  "00000110111110";
		Trees_din <= x"0bfe8f04";
		wait for Clk_period;
		Addr <=  "00000110111111";
		Trees_din <= x"ffa50715";
		wait for Clk_period;
		Addr <=  "00000111000000";
		Trees_din <= x"fff50715";
		wait for Clk_period;
		Addr <=  "00000111000001";
		Trees_din <= x"08005904";
		wait for Clk_period;
		Addr <=  "00000111000010";
		Trees_din <= x"00a30715";
		wait for Clk_period;
		Addr <=  "00000111000011";
		Trees_din <= x"00110715";
		wait for Clk_period;
		Addr <=  "00000111000100";
		Trees_din <= x"00250715";
		wait for Clk_period;
		Addr <=  "00000111000101";
		Trees_din <= x"000b0b2c";
		wait for Clk_period;
		Addr <=  "00000111000110";
		Trees_din <= x"00054904";
		wait for Clk_period;
		Addr <=  "00000111000111";
		Trees_din <= x"ff6607f1";
		wait for Clk_period;
		Addr <=  "00000111001000";
		Trees_din <= x"03ff4c1c";
		wait for Clk_period;
		Addr <=  "00000111001001";
		Trees_din <= x"15048510";
		wait for Clk_period;
		Addr <=  "00000111001010";
		Trees_din <= x"08005408";
		wait for Clk_period;
		Addr <=  "00000111001011";
		Trees_din <= x"07004e04";
		wait for Clk_period;
		Addr <=  "00000111001100";
		Trees_din <= x"ffea07f1";
		wait for Clk_period;
		Addr <=  "00000111001101";
		Trees_din <= x"ff5d07f1";
		wait for Clk_period;
		Addr <=  "00000111001110";
		Trees_din <= x"000a0704";
		wait for Clk_period;
		Addr <=  "00000111001111";
		Trees_din <= x"ff8c07f1";
		wait for Clk_period;
		Addr <=  "00000111010000";
		Trees_din <= x"002a07f1";
		wait for Clk_period;
		Addr <=  "00000111010001";
		Trees_din <= x"04fedf04";
		wait for Clk_period;
		Addr <=  "00000111010010";
		Trees_din <= x"ff9307f1";
		wait for Clk_period;
		Addr <=  "00000111010011";
		Trees_din <= x"08005204";
		wait for Clk_period;
		Addr <=  "00000111010100";
		Trees_din <= x"00a907f1";
		wait for Clk_period;
		Addr <=  "00000111010101";
		Trees_din <= x"001207f1";
		wait for Clk_period;
		Addr <=  "00000111010110";
		Trees_din <= x"1f040004";
		wait for Clk_period;
		Addr <=  "00000111010111";
		Trees_din <= x"ffe407f1";
		wait for Clk_period;
		Addr <=  "00000111011000";
		Trees_din <= x"0f024c04";
		wait for Clk_period;
		Addr <=  "00000111011001";
		Trees_din <= x"008307f1";
		wait for Clk_period;
		Addr <=  "00000111011010";
		Trees_din <= x"001907f1";
		wait for Clk_period;
		Addr <=  "00000111011011";
		Trees_din <= x"000e0630";
		wait for Clk_period;
		Addr <=  "00000111011100";
		Trees_din <= x"03fd461c";
		wait for Clk_period;
		Addr <=  "00000111011101";
		Trees_din <= x"0904f30c";
		wait for Clk_period;
		Addr <=  "00000111011110";
		Trees_din <= x"03fd3608";
		wait for Clk_period;
		Addr <=  "00000111011111";
		Trees_din <= x"02feff04";
		wait for Clk_period;
		Addr <=  "00000111100000";
		Trees_din <= x"ffe307f1";
		wait for Clk_period;
		Addr <=  "00000111100001";
		Trees_din <= x"008107f1";
		wait for Clk_period;
		Addr <=  "00000111100010";
		Trees_din <= x"ff8c07f1";
		wait for Clk_period;
		Addr <=  "00000111100011";
		Trees_din <= x"05072408";
		wait for Clk_period;
		Addr <=  "00000111100100";
		Trees_din <= x"14036304";
		wait for Clk_period;
		Addr <=  "00000111100101";
		Trees_din <= x"006c07f1";
		wait for Clk_period;
		Addr <=  "00000111100110";
		Trees_din <= x"fff907f1";
		wait for Clk_period;
		Addr <=  "00000111100111";
		Trees_din <= x"0c00da04";
		wait for Clk_period;
		Addr <=  "00000111101000";
		Trees_din <= x"ff5b07f1";
		wait for Clk_period;
		Addr <=  "00000111101001";
		Trees_din <= x"ffdd07f1";
		wait for Clk_period;
		Addr <=  "00000111101010";
		Trees_din <= x"0d001104";
		wait for Clk_period;
		Addr <=  "00000111101011";
		Trees_din <= x"fff507f1";
		wait for Clk_period;
		Addr <=  "00000111101100";
		Trees_din <= x"0b041c08";
		wait for Clk_period;
		Addr <=  "00000111101101";
		Trees_din <= x"1b03dd04";
		wait for Clk_period;
		Addr <=  "00000111101110";
		Trees_din <= x"00a107f1";
		wait for Clk_period;
		Addr <=  "00000111101111";
		Trees_din <= x"000807f1";
		wait for Clk_period;
		Addr <=  "00000111110000";
		Trees_din <= x"10034504";
		wait for Clk_period;
		Addr <=  "00000111110001";
		Trees_din <= x"005b07f1";
		wait for Clk_period;
		Addr <=  "00000111110010";
		Trees_din <= x"ffbd07f1";
		wait for Clk_period;
		Addr <=  "00000111110011";
		Trees_din <= x"04078910";
		wait for Clk_period;
		Addr <=  "00000111110100";
		Trees_din <= x"0508d704";
		wait for Clk_period;
		Addr <=  "00000111110101";
		Trees_din <= x"00a507f1";
		wait for Clk_period;
		Addr <=  "00000111110110";
		Trees_din <= x"1a005508";
		wait for Clk_period;
		Addr <=  "00000111110111";
		Trees_din <= x"08005904";
		wait for Clk_period;
		Addr <=  "00000111111000";
		Trees_din <= x"009c07f1";
		wait for Clk_period;
		Addr <=  "00000111111001";
		Trees_din <= x"fff607f1";
		wait for Clk_period;
		Addr <=  "00000111111010";
		Trees_din <= x"ffa507f1";
		wait for Clk_period;
		Addr <=  "00000111111011";
		Trees_din <= x"001f07f1";
		wait for Clk_period;
		Addr <=  "00000111111100";
		Trees_din <= x"000b0b1c";
		wait for Clk_period;
		Addr <=  "00000111111101";
		Trees_din <= x"00054904";
		wait for Clk_period;
		Addr <=  "00000111111110";
		Trees_din <= x"ff6808a5";
		wait for Clk_period;
		Addr <=  "00000111111111";
		Trees_din <= x"04fda904";
		wait for Clk_period;
		Addr <=  "00001000000000";
		Trees_din <= x"ff7a08a5";
		wait for Clk_period;
		Addr <=  "00001000000001";
		Trees_din <= x"0f02af0c";
		wait for Clk_period;
		Addr <=  "00001000000010";
		Trees_din <= x"03fc0304";
		wait for Clk_period;
		Addr <=  "00001000000011";
		Trees_din <= x"ffa708a5";
		wait for Clk_period;
		Addr <=  "00001000000100";
		Trees_din <= x"01f9f904";
		wait for Clk_period;
		Addr <=  "00001000000101";
		Trees_din <= x"ffec08a5";
		wait for Clk_period;
		Addr <=  "00001000000110";
		Trees_din <= x"006c08a5";
		wait for Clk_period;
		Addr <=  "00001000000111";
		Trees_din <= x"14036804";
		wait for Clk_period;
		Addr <=  "00001000001000";
		Trees_din <= x"ff6008a5";
		wait for Clk_period;
		Addr <=  "00001000001001";
		Trees_din <= x"002b08a5";
		wait for Clk_period;
		Addr <=  "00001000001010";
		Trees_din <= x"000e062c";
		wait for Clk_period;
		Addr <=  "00001000001011";
		Trees_din <= x"03fddd20";
		wait for Clk_period;
		Addr <=  "00001000001100";
		Trees_din <= x"0a013710";
		wait for Clk_period;
		Addr <=  "00001000001101";
		Trees_din <= x"0a001408";
		wait for Clk_period;
		Addr <=  "00001000001110";
		Trees_din <= x"08005704";
		wait for Clk_period;
		Addr <=  "00001000001111";
		Trees_din <= x"004708a5";
		wait for Clk_period;
		Addr <=  "00001000010000";
		Trees_din <= x"ff6b08a5";
		wait for Clk_period;
		Addr <=  "00001000010001";
		Trees_din <= x"09054304";
		wait for Clk_period;
		Addr <=  "00001000010010";
		Trees_din <= x"00b808a5";
		wait for Clk_period;
		Addr <=  "00001000010011";
		Trees_din <= x"fffc08a5";
		wait for Clk_period;
		Addr <=  "00001000010100";
		Trees_din <= x"12009608";
		wait for Clk_period;
		Addr <=  "00001000010101";
		Trees_din <= x"07005404";
		wait for Clk_period;
		Addr <=  "00001000010110";
		Trees_din <= x"ff3408a5";
		wait for Clk_period;
		Addr <=  "00001000010111";
		Trees_din <= x"001908a5";
		wait for Clk_period;
		Addr <=  "00001000011000";
		Trees_din <= x"0a01f104";
		wait for Clk_period;
		Addr <=  "00001000011001";
		Trees_din <= x"ffda08a5";
		wait for Clk_period;
		Addr <=  "00001000011010";
		Trees_din <= x"006e08a5";
		wait for Clk_period;
		Addr <=  "00001000011011";
		Trees_din <= x"04fd5b08";
		wait for Clk_period;
		Addr <=  "00001000011100";
		Trees_din <= x"0b022604";
		wait for Clk_period;
		Addr <=  "00001000011101";
		Trees_din <= x"006808a5";
		wait for Clk_period;
		Addr <=  "00001000011110";
		Trees_din <= x"ff9c08a5";
		wait for Clk_period;
		Addr <=  "00001000011111";
		Trees_din <= x"009f08a5";
		wait for Clk_period;
		Addr <=  "00001000100000";
		Trees_din <= x"0508d708";
		wait for Clk_period;
		Addr <=  "00001000100001";
		Trees_din <= x"04078904";
		wait for Clk_period;
		Addr <=  "00001000100010";
		Trees_din <= x"00a208a5";
		wait for Clk_period;
		Addr <=  "00001000100011";
		Trees_din <= x"001d08a5";
		wait for Clk_period;
		Addr <=  "00001000100100";
		Trees_din <= x"1d009304";
		wait for Clk_period;
		Addr <=  "00001000100101";
		Trees_din <= x"ffbf08a5";
		wait for Clk_period;
		Addr <=  "00001000100110";
		Trees_din <= x"0b03b504";
		wait for Clk_period;
		Addr <=  "00001000100111";
		Trees_din <= x"009508a5";
		wait for Clk_period;
		Addr <=  "00001000101000";
		Trees_din <= x"000608a5";
		wait for Clk_period;
		Addr <=  "00001000101001";
		Trees_din <= x"000b0b28";
		wait for Clk_period;
		Addr <=  "00001000101010";
		Trees_din <= x"00054904";
		wait for Clk_period;
		Addr <=  "00001000101011";
		Trees_din <= x"ff690969";
		wait for Clk_period;
		Addr <=  "00001000101100";
		Trees_din <= x"04fda904";
		wait for Clk_period;
		Addr <=  "00001000101101";
		Trees_din <= x"ff800969";
		wait for Clk_period;
		Addr <=  "00001000101110";
		Trees_din <= x"01fb6610";
		wait for Clk_period;
		Addr <=  "00001000101111";
		Trees_din <= x"1e006408";
		wait for Clk_period;
		Addr <=  "00001000110000";
		Trees_din <= x"09046104";
		wait for Clk_period;
		Addr <=  "00001000110001";
		Trees_din <= x"001d0969";
		wait for Clk_period;
		Addr <=  "00001000110010";
		Trees_din <= x"009b0969";
		wait for Clk_period;
		Addr <=  "00001000110011";
		Trees_din <= x"17004704";
		wait for Clk_period;
		Addr <=  "00001000110100";
		Trees_din <= x"ff960969";
		wait for Clk_period;
		Addr <=  "00001000110101";
		Trees_din <= x"00380969";
		wait for Clk_period;
		Addr <=  "00001000110110";
		Trees_din <= x"1c003508";
		wait for Clk_period;
		Addr <=  "00001000110111";
		Trees_din <= x"1100ef04";
		wait for Clk_period;
		Addr <=  "00001000111000";
		Trees_din <= x"ffde0969";
		wait for Clk_period;
		Addr <=  "00001000111001";
		Trees_din <= x"ff6e0969";
		wait for Clk_period;
		Addr <=  "00001000111010";
		Trees_din <= x"03fd0f04";
		wait for Clk_period;
		Addr <=  "00001000111011";
		Trees_din <= x"ffc90969";
		wait for Clk_period;
		Addr <=  "00001000111100";
		Trees_din <= x"00590969";
		wait for Clk_period;
		Addr <=  "00001000111101";
		Trees_din <= x"000ec830";
		wait for Clk_period;
		Addr <=  "00001000111110";
		Trees_din <= x"03fd461c";
		wait for Clk_period;
		Addr <=  "00001000111111";
		Trees_din <= x"01fcd510";
		wait for Clk_period;
		Addr <=  "00001001000000";
		Trees_din <= x"08005108";
		wait for Clk_period;
		Addr <=  "00001001000001";
		Trees_din <= x"1c002304";
		wait for Clk_period;
		Addr <=  "00001001000010";
		Trees_din <= x"000f0969";
		wait for Clk_period;
		Addr <=  "00001001000011";
		Trees_din <= x"00860969";
		wait for Clk_period;
		Addr <=  "00001001000100";
		Trees_din <= x"06fd7204";
		wait for Clk_period;
		Addr <=  "00001001000101";
		Trees_din <= x"00130969";
		wait for Clk_period;
		Addr <=  "00001001000110";
		Trees_din <= x"ff740969";
		wait for Clk_period;
		Addr <=  "00001001000111";
		Trees_din <= x"03fac204";
		wait for Clk_period;
		Addr <=  "00001001001000";
		Trees_din <= x"fff60969";
		wait for Clk_period;
		Addr <=  "00001001001001";
		Trees_din <= x"07005c04";
		wait for Clk_period;
		Addr <=  "00001001001010";
		Trees_din <= x"00980969";
		wait for Clk_period;
		Addr <=  "00001001001011";
		Trees_din <= x"002a0969";
		wait for Clk_period;
		Addr <=  "00001001001100";
		Trees_din <= x"06fc9b10";
		wait for Clk_period;
		Addr <=  "00001001001101";
		Trees_din <= x"1b024108";
		wait for Clk_period;
		Addr <=  "00001001001110";
		Trees_din <= x"0a000304";
		wait for Clk_period;
		Addr <=  "00001001001111";
		Trees_din <= x"ffff0969";
		wait for Clk_period;
		Addr <=  "00001001010000";
		Trees_din <= x"00910969";
		wait for Clk_period;
		Addr <=  "00001001010001";
		Trees_din <= x"02fed204";
		wait for Clk_period;
		Addr <=  "00001001010010";
		Trees_din <= x"ff740969";
		wait for Clk_period;
		Addr <=  "00001001010011";
		Trees_din <= x"00540969";
		wait for Clk_period;
		Addr <=  "00001001010100";
		Trees_din <= x"009b0969";
		wait for Clk_period;
		Addr <=  "00001001010101";
		Trees_din <= x"03fafa04";
		wait for Clk_period;
		Addr <=  "00001001010110";
		Trees_din <= x"00040969";
		wait for Clk_period;
		Addr <=  "00001001010111";
		Trees_din <= x"04078904";
		wait for Clk_period;
		Addr <=  "00001001011000";
		Trees_din <= x"00a00969";
		wait for Clk_period;
		Addr <=  "00001001011001";
		Trees_din <= x"00050969";
		wait for Clk_period;
		Addr <=  "00001001011010";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00001001011011";
		Trees_din <= x"000b0b28";
		wait for Clk_period;
		Addr <=  "00001001011100";
		Trees_din <= x"00054904";
		wait for Clk_period;
		Addr <=  "00001001011101";
		Trees_din <= x"ff6b0a31";
		wait for Clk_period;
		Addr <=  "00001001011110";
		Trees_din <= x"03ff4c18";
		wait for Clk_period;
		Addr <=  "00001001011111";
		Trees_din <= x"15048510";
		wait for Clk_period;
		Addr <=  "00001001100000";
		Trees_din <= x"08005608";
		wait for Clk_period;
		Addr <=  "00001001100001";
		Trees_din <= x"0c028704";
		wait for Clk_period;
		Addr <=  "00001001100010";
		Trees_din <= x"ff670a31";
		wait for Clk_period;
		Addr <=  "00001001100011";
		Trees_din <= x"fff10a31";
		wait for Clk_period;
		Addr <=  "00001001100100";
		Trees_din <= x"00097504";
		wait for Clk_period;
		Addr <=  "00001001100101";
		Trees_din <= x"ff9e0a31";
		wait for Clk_period;
		Addr <=  "00001001100110";
		Trees_din <= x"00220a31";
		wait for Clk_period;
		Addr <=  "00001001100111";
		Trees_din <= x"04fedf04";
		wait for Clk_period;
		Addr <=  "00001001101000";
		Trees_din <= x"ffa90a31";
		wait for Clk_period;
		Addr <=  "00001001101001";
		Trees_din <= x"00640a31";
		wait for Clk_period;
		Addr <=  "00001001101010";
		Trees_din <= x"1b014408";
		wait for Clk_period;
		Addr <=  "00001001101011";
		Trees_din <= x"11005304";
		wait for Clk_period;
		Addr <=  "00001001101100";
		Trees_din <= x"004e0a31";
		wait for Clk_period;
		Addr <=  "00001001101101";
		Trees_din <= x"ffa70a31";
		wait for Clk_period;
		Addr <=  "00001001101110";
		Trees_din <= x"00670a31";
		wait for Clk_period;
		Addr <=  "00001001101111";
		Trees_din <= x"000ec830";
		wait for Clk_period;
		Addr <=  "00001001110000";
		Trees_din <= x"03fd461c";
		wait for Clk_period;
		Addr <=  "00001001110001";
		Trees_din <= x"01fcd510";
		wait for Clk_period;
		Addr <=  "00001001110010";
		Trees_din <= x"08005108";
		wait for Clk_period;
		Addr <=  "00001001110011";
		Trees_din <= x"1c002304";
		wait for Clk_period;
		Addr <=  "00001001110100";
		Trees_din <= x"000e0a31";
		wait for Clk_period;
		Addr <=  "00001001110101";
		Trees_din <= x"00790a31";
		wait for Clk_period;
		Addr <=  "00001001110110";
		Trees_din <= x"11003904";
		wait for Clk_period;
		Addr <=  "00001001110111";
		Trees_din <= x"ff4f0a31";
		wait for Clk_period;
		Addr <=  "00001001111000";
		Trees_din <= x"fff60a31";
		wait for Clk_period;
		Addr <=  "00001001111001";
		Trees_din <= x"03fac204";
		wait for Clk_period;
		Addr <=  "00001001111010";
		Trees_din <= x"fff60a31";
		wait for Clk_period;
		Addr <=  "00001001111011";
		Trees_din <= x"09051d04";
		wait for Clk_period;
		Addr <=  "00001001111100";
		Trees_din <= x"00910a31";
		wait for Clk_period;
		Addr <=  "00001001111101";
		Trees_din <= x"001c0a31";
		wait for Clk_period;
		Addr <=  "00001001111110";
		Trees_din <= x"06fc9b10";
		wait for Clk_period;
		Addr <=  "00001001111111";
		Trees_din <= x"19009308";
		wait for Clk_period;
		Addr <=  "00001010000000";
		Trees_din <= x"19008e04";
		wait for Clk_period;
		Addr <=  "00001010000001";
		Trees_din <= x"00560a31";
		wait for Clk_period;
		Addr <=  "00001010000010";
		Trees_din <= x"ff6d0a31";
		wait for Clk_period;
		Addr <=  "00001010000011";
		Trees_din <= x"15047004";
		wait for Clk_period;
		Addr <=  "00001010000100";
		Trees_din <= x"00860a31";
		wait for Clk_period;
		Addr <=  "00001010000101";
		Trees_din <= x"001b0a31";
		wait for Clk_period;
		Addr <=  "00001010000110";
		Trees_din <= x"00960a31";
		wait for Clk_period;
		Addr <=  "00001010000111";
		Trees_din <= x"03fafa04";
		wait for Clk_period;
		Addr <=  "00001010001000";
		Trees_din <= x"00000a31";
		wait for Clk_period;
		Addr <=  "00001010001001";
		Trees_din <= x"04078904";
		wait for Clk_period;
		Addr <=  "00001010001010";
		Trees_din <= x"009e0a31";
		wait for Clk_period;
		Addr <=  "00001010001011";
		Trees_din <= x"00020a31";
		wait for Clk_period;
		Addr <=  "00001010001100";
		Trees_din <= x"000bb830";
		wait for Clk_period;
		Addr <=  "00001010001101";
		Trees_din <= x"00054904";
		wait for Clk_period;
		Addr <=  "00001010001110";
		Trees_din <= x"ff6c0aed";
		wait for Clk_period;
		Addr <=  "00001010001111";
		Trees_din <= x"04fee81c";
		wait for Clk_period;
		Addr <=  "00001010010000";
		Trees_din <= x"1000ae10";
		wait for Clk_period;
		Addr <=  "00001010010001";
		Trees_din <= x"01fa3b08";
		wait for Clk_period;
		Addr <=  "00001010010010";
		Trees_din <= x"1b030204";
		wait for Clk_period;
		Addr <=  "00001010010011";
		Trees_din <= x"00050aed";
		wait for Clk_period;
		Addr <=  "00001010010100";
		Trees_din <= x"005b0aed";
		wait for Clk_period;
		Addr <=  "00001010010101";
		Trees_din <= x"0bfe4804";
		wait for Clk_period;
		Addr <=  "00001010010110";
		Trees_din <= x"ffa40aed";
		wait for Clk_period;
		Addr <=  "00001010010111";
		Trees_din <= x"fff90aed";
		wait for Clk_period;
		Addr <=  "00001010011000";
		Trees_din <= x"1900a708";
		wait for Clk_period;
		Addr <=  "00001010011001";
		Trees_din <= x"1a004204";
		wait for Clk_period;
		Addr <=  "00001010011010";
		Trees_din <= x"ffcd0aed";
		wait for Clk_period;
		Addr <=  "00001010011011";
		Trees_din <= x"ff6a0aed";
		wait for Clk_period;
		Addr <=  "00001010011100";
		Trees_din <= x"00100aed";
		wait for Clk_period;
		Addr <=  "00001010011101";
		Trees_din <= x"0b03f40c";
		wait for Clk_period;
		Addr <=  "00001010011110";
		Trees_din <= x"05fb7b04";
		wait for Clk_period;
		Addr <=  "00001010011111";
		Trees_din <= x"ffcf0aed";
		wait for Clk_period;
		Addr <=  "00001010100000";
		Trees_din <= x"06fe5504";
		wait for Clk_period;
		Addr <=  "00001010100001";
		Trees_din <= x"007a0aed";
		wait for Clk_period;
		Addr <=  "00001010100010";
		Trees_din <= x"fff80aed";
		wait for Clk_period;
		Addr <=  "00001010100011";
		Trees_din <= x"ffa70aed";
		wait for Clk_period;
		Addr <=  "00001010100100";
		Trees_din <= x"000ec824";
		wait for Clk_period;
		Addr <=  "00001010100101";
		Trees_din <= x"02faa208";
		wait for Clk_period;
		Addr <=  "00001010100110";
		Trees_din <= x"02fa2c04";
		wait for Clk_period;
		Addr <=  "00001010100111";
		Trees_din <= x"00590aed";
		wait for Clk_period;
		Addr <=  "00001010101000";
		Trees_din <= x"ff440aed";
		wait for Clk_period;
		Addr <=  "00001010101001";
		Trees_din <= x"03fbf710";
		wait for Clk_period;
		Addr <=  "00001010101010";
		Trees_din <= x"01fbc708";
		wait for Clk_period;
		Addr <=  "00001010101011";
		Trees_din <= x"19008f04";
		wait for Clk_period;
		Addr <=  "00001010101100";
		Trees_din <= x"ff220aed";
		wait for Clk_period;
		Addr <=  "00001010101101";
		Trees_din <= x"00230aed";
		wait for Clk_period;
		Addr <=  "00001010101110";
		Trees_din <= x"15fa8d04";
		wait for Clk_period;
		Addr <=  "00001010101111";
		Trees_din <= x"00050aed";
		wait for Clk_period;
		Addr <=  "00001010110000";
		Trees_din <= x"00710aed";
		wait for Clk_period;
		Addr <=  "00001010110001";
		Trees_din <= x"08005c08";
		wait for Clk_period;
		Addr <=  "00001010110010";
		Trees_din <= x"1504f204";
		wait for Clk_period;
		Addr <=  "00001010110011";
		Trees_din <= x"008f0aed";
		wait for Clk_period;
		Addr <=  "00001010110100";
		Trees_din <= x"001c0aed";
		wait for Clk_period;
		Addr <=  "00001010110101";
		Trees_din <= x"ffb90aed";
		wait for Clk_period;
		Addr <=  "00001010110110";
		Trees_din <= x"03fafa04";
		wait for Clk_period;
		Addr <=  "00001010110111";
		Trees_din <= x"fffd0aed";
		wait for Clk_period;
		Addr <=  "00001010111000";
		Trees_din <= x"04078904";
		wait for Clk_period;
		Addr <=  "00001010111001";
		Trees_din <= x"009d0aed";
		wait for Clk_period;
		Addr <=  "00001010111010";
		Trees_din <= x"00010aed";
		wait for Clk_period;
		Addr <=  "00001010111011";
		Trees_din <= x"000c1020";
		wait for Clk_period;
		Addr <=  "00001010111100";
		Trees_din <= x"00054904";
		wait for Clk_period;
		Addr <=  "00001010111101";
		Trees_din <= x"ff6e0b79";
		wait for Clk_period;
		Addr <=  "00001010111110";
		Trees_din <= x"06fa6a04";
		wait for Clk_period;
		Addr <=  "00001010111111";
		Trees_din <= x"00600b79";
		wait for Clk_period;
		Addr <=  "00001011000000";
		Trees_din <= x"03000310";
		wait for Clk_period;
		Addr <=  "00001011000001";
		Trees_din <= x"15057c08";
		wait for Clk_period;
		Addr <=  "00001011000010";
		Trees_din <= x"08004c04";
		wait for Clk_period;
		Addr <=  "00001011000011";
		Trees_din <= x"00150b79";
		wait for Clk_period;
		Addr <=  "00001011000100";
		Trees_din <= x"ffb40b79";
		wait for Clk_period;
		Addr <=  "00001011000101";
		Trees_din <= x"0c00bc04";
		wait for Clk_period;
		Addr <=  "00001011000110";
		Trees_din <= x"00690b79";
		wait for Clk_period;
		Addr <=  "00001011000111";
		Trees_din <= x"fff10b79";
		wait for Clk_period;
		Addr <=  "00001011001000";
		Trees_din <= x"09041004";
		wait for Clk_period;
		Addr <=  "00001011001001";
		Trees_din <= x"005f0b79";
		wait for Clk_period;
		Addr <=  "00001011001010";
		Trees_din <= x"fff80b79";
		wait for Clk_period;
		Addr <=  "00001011001011";
		Trees_din <= x"000ec81c";
		wait for Clk_period;
		Addr <=  "00001011001100";
		Trees_din <= x"02faa208";
		wait for Clk_period;
		Addr <=  "00001011001101";
		Trees_din <= x"02fa1704";
		wait for Clk_period;
		Addr <=  "00001011001110";
		Trees_din <= x"00630b79";
		wait for Clk_period;
		Addr <=  "00001011001111";
		Trees_din <= x"ff610b79";
		wait for Clk_period;
		Addr <=  "00001011010000";
		Trees_din <= x"03fd4610";
		wait for Clk_period;
		Addr <=  "00001011010001";
		Trees_din <= x"0d01f708";
		wait for Clk_period;
		Addr <=  "00001011010010";
		Trees_din <= x"0904a904";
		wait for Clk_period;
		Addr <=  "00001011010011";
		Trees_din <= x"008a0b79";
		wait for Clk_period;
		Addr <=  "00001011010100";
		Trees_din <= x"001b0b79";
		wait for Clk_period;
		Addr <=  "00001011010101";
		Trees_din <= x"17004204";
		wait for Clk_period;
		Addr <=  "00001011010110";
		Trees_din <= x"00400b79";
		wait for Clk_period;
		Addr <=  "00001011010111";
		Trees_din <= x"ff9f0b79";
		wait for Clk_period;
		Addr <=  "00001011011000";
		Trees_din <= x"00900b79";
		wait for Clk_period;
		Addr <=  "00001011011001";
		Trees_din <= x"03fafa04";
		wait for Clk_period;
		Addr <=  "00001011011010";
		Trees_din <= x"fffd0b79";
		wait for Clk_period;
		Addr <=  "00001011011011";
		Trees_din <= x"04078904";
		wait for Clk_period;
		Addr <=  "00001011011100";
		Trees_din <= x"009b0b79";
		wait for Clk_period;
		Addr <=  "00001011011101";
		Trees_din <= x"00000b79";
		wait for Clk_period;
		Addr <=  "00001011011110";
		Trees_din <= x"000c1030";
		wait for Clk_period;
		Addr <=  "00001011011111";
		Trees_din <= x"00071308";
		wait for Clk_period;
		Addr <=  "00001011100000";
		Trees_din <= x"1900af04";
		wait for Clk_period;
		Addr <=  "00001011100001";
		Trees_din <= x"ff740c35";
		wait for Clk_period;
		Addr <=  "00001011100010";
		Trees_din <= x"ffdf0c35";
		wait for Clk_period;
		Addr <=  "00001011100011";
		Trees_din <= x"04fee814";
		wait for Clk_period;
		Addr <=  "00001011100100";
		Trees_din <= x"1c00370c";
		wait for Clk_period;
		Addr <=  "00001011100101";
		Trees_din <= x"18003a08";
		wait for Clk_period;
		Addr <=  "00001011100110";
		Trees_din <= x"08005504";
		wait for Clk_period;
		Addr <=  "00001011100111";
		Trees_din <= x"ffbf0c35";
		wait for Clk_period;
		Addr <=  "00001011101000";
		Trees_din <= x"001e0c35";
		wait for Clk_period;
		Addr <=  "00001011101001";
		Trees_din <= x"00590c35";
		wait for Clk_period;
		Addr <=  "00001011101010";
		Trees_din <= x"10000f04";
		wait for Clk_period;
		Addr <=  "00001011101011";
		Trees_din <= x"00000c35";
		wait for Clk_period;
		Addr <=  "00001011101100";
		Trees_din <= x"ff6d0c35";
		wait for Clk_period;
		Addr <=  "00001011101101";
		Trees_din <= x"06ff180c";
		wait for Clk_period;
		Addr <=  "00001011101110";
		Trees_din <= x"1d00ad04";
		wait for Clk_period;
		Addr <=  "00001011101111";
		Trees_din <= x"ffe80c35";
		wait for Clk_period;
		Addr <=  "00001011110000";
		Trees_din <= x"05fe2a04";
		wait for Clk_period;
		Addr <=  "00001011110001";
		Trees_din <= x"00100c35";
		wait for Clk_period;
		Addr <=  "00001011110010";
		Trees_din <= x"007e0c35";
		wait for Clk_period;
		Addr <=  "00001011110011";
		Trees_din <= x"0e016504";
		wait for Clk_period;
		Addr <=  "00001011110100";
		Trees_din <= x"00210c35";
		wait for Clk_period;
		Addr <=  "00001011110101";
		Trees_din <= x"ff860c35";
		wait for Clk_period;
		Addr <=  "00001011110110";
		Trees_din <= x"000ec820";
		wait for Clk_period;
		Addr <=  "00001011110111";
		Trees_din <= x"02faa208";
		wait for Clk_period;
		Addr <=  "00001011111000";
		Trees_din <= x"02fa2c04";
		wait for Clk_period;
		Addr <=  "00001011111001";
		Trees_din <= x"004c0c35";
		wait for Clk_period;
		Addr <=  "00001011111010";
		Trees_din <= x"ff590c35";
		wait for Clk_period;
		Addr <=  "00001011111011";
		Trees_din <= x"03fc920c";
		wait for Clk_period;
		Addr <=  "00001011111100";
		Trees_din <= x"01fc3108";
		wait for Clk_period;
		Addr <=  "00001011111101";
		Trees_din <= x"06fcef04";
		wait for Clk_period;
		Addr <=  "00001011111110";
		Trees_din <= x"002f0c35";
		wait for Clk_period;
		Addr <=  "00001011111111";
		Trees_din <= x"ff6c0c35";
		wait for Clk_period;
		Addr <=  "00001100000000";
		Trees_din <= x"006d0c35";
		wait for Clk_period;
		Addr <=  "00001100000001";
		Trees_din <= x"09f76208";
		wait for Clk_period;
		Addr <=  "00001100000010";
		Trees_din <= x"1302e204";
		wait for Clk_period;
		Addr <=  "00001100000011";
		Trees_din <= x"00540c35";
		wait for Clk_period;
		Addr <=  "00001100000100";
		Trees_din <= x"ffb20c35";
		wait for Clk_period;
		Addr <=  "00001100000101";
		Trees_din <= x"008f0c35";
		wait for Clk_period;
		Addr <=  "00001100000110";
		Trees_din <= x"0c03ed0c";
		wait for Clk_period;
		Addr <=  "00001100000111";
		Trees_din <= x"09f71e08";
		wait for Clk_period;
		Addr <=  "00001100001000";
		Trees_din <= x"12009204";
		wait for Clk_period;
		Addr <=  "00001100001001";
		Trees_din <= x"fffb0c35";
		wait for Clk_period;
		Addr <=  "00001100001010";
		Trees_din <= x"00550c35";
		wait for Clk_period;
		Addr <=  "00001100001011";
		Trees_din <= x"009b0c35";
		wait for Clk_period;
		Addr <=  "00001100001100";
		Trees_din <= x"000f0c35";
		wait for Clk_period;
		Addr <=  "00001100001101";
		Trees_din <= x"000c1020";
		wait for Clk_period;
		Addr <=  "00001100001110";
		Trees_din <= x"00054904";
		wait for Clk_period;
		Addr <=  "00001100001111";
		Trees_din <= x"ff730cd1";
		wait for Clk_period;
		Addr <=  "00001100010000";
		Trees_din <= x"06fa6a04";
		wait for Clk_period;
		Addr <=  "00001100010001";
		Trees_din <= x"00560cd1";
		wait for Clk_period;
		Addr <=  "00001100010010";
		Trees_din <= x"03fdfa0c";
		wait for Clk_period;
		Addr <=  "00001100010011";
		Trees_din <= x"15057c08";
		wait for Clk_period;
		Addr <=  "00001100010100";
		Trees_din <= x"08005604";
		wait for Clk_period;
		Addr <=  "00001100010101";
		Trees_din <= x"ff960cd1";
		wait for Clk_period;
		Addr <=  "00001100010110";
		Trees_din <= x"fff10cd1";
		wait for Clk_period;
		Addr <=  "00001100010111";
		Trees_din <= x"003d0cd1";
		wait for Clk_period;
		Addr <=  "00001100011000";
		Trees_din <= x"0c014d08";
		wait for Clk_period;
		Addr <=  "00001100011001";
		Trees_din <= x"18004004";
		wait for Clk_period;
		Addr <=  "00001100011010";
		Trees_din <= x"ffb50cd1";
		wait for Clk_period;
		Addr <=  "00001100011011";
		Trees_din <= x"00290cd1";
		wait for Clk_period;
		Addr <=  "00001100011100";
		Trees_din <= x"00540cd1";
		wait for Clk_period;
		Addr <=  "00001100011101";
		Trees_din <= x"000ec824";
		wait for Clk_period;
		Addr <=  "00001100011110";
		Trees_din <= x"0d01fb10";
		wait for Clk_period;
		Addr <=  "00001100011111";
		Trees_din <= x"050c4e08";
		wait for Clk_period;
		Addr <=  "00001100100000";
		Trees_din <= x"15f96b04";
		wait for Clk_period;
		Addr <=  "00001100100001";
		Trees_din <= x"00280cd1";
		wait for Clk_period;
		Addr <=  "00001100100010";
		Trees_din <= x"008f0cd1";
		wait for Clk_period;
		Addr <=  "00001100100011";
		Trees_din <= x"09039e04";
		wait for Clk_period;
		Addr <=  "00001100100100";
		Trees_din <= x"005c0cd1";
		wait for Clk_period;
		Addr <=  "00001100100101";
		Trees_din <= x"ffaf0cd1";
		wait for Clk_period;
		Addr <=  "00001100100110";
		Trees_din <= x"1200980c";
		wait for Clk_period;
		Addr <=  "00001100100111";
		Trees_din <= x"08005304";
		wait for Clk_period;
		Addr <=  "00001100101000";
		Trees_din <= x"ff1a0cd1";
		wait for Clk_period;
		Addr <=  "00001100101001";
		Trees_din <= x"05081c04";
		wait for Clk_period;
		Addr <=  "00001100101010";
		Trees_din <= x"00450cd1";
		wait for Clk_period;
		Addr <=  "00001100101011";
		Trees_din <= x"ffc40cd1";
		wait for Clk_period;
		Addr <=  "00001100101100";
		Trees_din <= x"14017e04";
		wait for Clk_period;
		Addr <=  "00001100101101";
		Trees_din <= x"00770cd1";
		wait for Clk_period;
		Addr <=  "00001100101110";
		Trees_din <= x"fffc0cd1";
		wait for Clk_period;
		Addr <=  "00001100101111";
		Trees_din <= x"0c03ed08";
		wait for Clk_period;
		Addr <=  "00001100110000";
		Trees_din <= x"09f71e04";
		wait for Clk_period;
		Addr <=  "00001100110001";
		Trees_din <= x"00300cd1";
		wait for Clk_period;
		Addr <=  "00001100110010";
		Trees_din <= x"009a0cd1";
		wait for Clk_period;
		Addr <=  "00001100110011";
		Trees_din <= x"000c0cd1";
		wait for Clk_period;
		Addr <=  "00001100110100";
		Trees_din <= x"000ec83c";
		wait for Clk_period;
		Addr <=  "00001100110101";
		Trees_din <= x"00087608";
		wait for Clk_period;
		Addr <=  "00001100110110";
		Trees_din <= x"15056004";
		wait for Clk_period;
		Addr <=  "00001100110111";
		Trees_din <= x"ff7f0d5d";
		wait for Clk_period;
		Addr <=  "00001100111000";
		Trees_din <= x"fff40d5d";
		wait for Clk_period;
		Addr <=  "00001100111001";
		Trees_din <= x"0a01371c";
		wait for Clk_period;
		Addr <=  "00001100111010";
		Trees_din <= x"0a001410";
		wait for Clk_period;
		Addr <=  "00001100111011";
		Trees_din <= x"0c00c508";
		wait for Clk_period;
		Addr <=  "00001100111100";
		Trees_din <= x"18003f04";
		wait for Clk_period;
		Addr <=  "00001100111101";
		Trees_din <= x"ff9d0d5d";
		wait for Clk_period;
		Addr <=  "00001100111110";
		Trees_din <= x"002d0d5d";
		wait for Clk_period;
		Addr <=  "00001100111111";
		Trees_din <= x"03fd2f04";
		wait for Clk_period;
		Addr <=  "00001101000000";
		Trees_din <= x"000d0d5d";
		wait for Clk_period;
		Addr <=  "00001101000001";
		Trees_din <= x"00530d5d";
		wait for Clk_period;
		Addr <=  "00001101000010";
		Trees_din <= x"0ffeb104";
		wait for Clk_period;
		Addr <=  "00001101000011";
		Trees_din <= x"00050d5d";
		wait for Clk_period;
		Addr <=  "00001101000100";
		Trees_din <= x"07005b04";
		wait for Clk_period;
		Addr <=  "00001101000101";
		Trees_din <= x"00830d5d";
		wait for Clk_period;
		Addr <=  "00001101000110";
		Trees_din <= x"00130d5d";
		wait for Clk_period;
		Addr <=  "00001101000111";
		Trees_din <= x"03fdea10";
		wait for Clk_period;
		Addr <=  "00001101001000";
		Trees_din <= x"10027808";
		wait for Clk_period;
		Addr <=  "00001101001001";
		Trees_din <= x"0a024804";
		wait for Clk_period;
		Addr <=  "00001101001010";
		Trees_din <= x"ffb90d5d";
		wait for Clk_period;
		Addr <=  "00001101001011";
		Trees_din <= x"004e0d5d";
		wait for Clk_period;
		Addr <=  "00001101001100";
		Trees_din <= x"12009d04";
		wait for Clk_period;
		Addr <=  "00001101001101";
		Trees_din <= x"ff5a0d5d";
		wait for Clk_period;
		Addr <=  "00001101001110";
		Trees_din <= x"002a0d5d";
		wait for Clk_period;
		Addr <=  "00001101001111";
		Trees_din <= x"14020a04";
		wait for Clk_period;
		Addr <=  "00001101010000";
		Trees_din <= x"00700d5d";
		wait for Clk_period;
		Addr <=  "00001101010001";
		Trees_din <= x"fffe0d5d";
		wait for Clk_period;
		Addr <=  "00001101010010";
		Trees_din <= x"0100fc08";
		wait for Clk_period;
		Addr <=  "00001101010011";
		Trees_din <= x"09f71e04";
		wait for Clk_period;
		Addr <=  "00001101010100";
		Trees_din <= x"00260d5d";
		wait for Clk_period;
		Addr <=  "00001101010101";
		Trees_din <= x"00990d5d";
		wait for Clk_period;
		Addr <=  "00001101010110";
		Trees_din <= x"00020d5d";
		wait for Clk_period;
		Addr <=  "00001101010111";
		Trees_din <= x"000ec834";
		wait for Clk_period;
		Addr <=  "00001101011000";
		Trees_din <= x"00054904";
		wait for Clk_period;
		Addr <=  "00001101011001";
		Trees_din <= x"ff7a0dd9";
		wait for Clk_period;
		Addr <=  "00001101011010";
		Trees_din <= x"03fde220";
		wait for Clk_period;
		Addr <=  "00001101011011";
		Trees_din <= x"0a013710";
		wait for Clk_period;
		Addr <=  "00001101011100";
		Trees_din <= x"0a001508";
		wait for Clk_period;
		Addr <=  "00001101011101";
		Trees_din <= x"0f016704";
		wait for Clk_period;
		Addr <=  "00001101011110";
		Trees_din <= x"ffba0dd9";
		wait for Clk_period;
		Addr <=  "00001101011111";
		Trees_din <= x"00250dd9";
		wait for Clk_period;
		Addr <=  "00001101100000";
		Trees_din <= x"000a8004";
		wait for Clk_period;
		Addr <=  "00001101100001";
		Trees_din <= x"ffd70dd9";
		wait for Clk_period;
		Addr <=  "00001101100010";
		Trees_din <= x"00650dd9";
		wait for Clk_period;
		Addr <=  "00001101100011";
		Trees_din <= x"0c00c208";
		wait for Clk_period;
		Addr <=  "00001101100100";
		Trees_din <= x"1c003f04";
		wait for Clk_period;
		Addr <=  "00001101100101";
		Trees_din <= x"00430dd9";
		wait for Clk_period;
		Addr <=  "00001101100110";
		Trees_din <= x"ffae0dd9";
		wait for Clk_period;
		Addr <=  "00001101100111";
		Trees_din <= x"08005404";
		wait for Clk_period;
		Addr <=  "00001101101000";
		Trees_din <= x"ff4b0dd9";
		wait for Clk_period;
		Addr <=  "00001101101001";
		Trees_din <= x"fffd0dd9";
		wait for Clk_period;
		Addr <=  "00001101101010";
		Trees_din <= x"000b0b08";
		wait for Clk_period;
		Addr <=  "00001101101011";
		Trees_din <= x"12009704";
		wait for Clk_period;
		Addr <=  "00001101101100";
		Trees_din <= x"00320dd9";
		wait for Clk_period;
		Addr <=  "00001101101101";
		Trees_din <= x"ffcd0dd9";
		wait for Clk_period;
		Addr <=  "00001101101110";
		Trees_din <= x"04fd5b04";
		wait for Clk_period;
		Addr <=  "00001101101111";
		Trees_din <= x"fff50dd9";
		wait for Clk_period;
		Addr <=  "00001101110000";
		Trees_din <= x"00820dd9";
		wait for Clk_period;
		Addr <=  "00001101110001";
		Trees_din <= x"05f92504";
		wait for Clk_period;
		Addr <=  "00001101110010";
		Trees_din <= x"00200dd9";
		wait for Clk_period;
		Addr <=  "00001101110011";
		Trees_din <= x"09f71e04";
		wait for Clk_period;
		Addr <=  "00001101110100";
		Trees_din <= x"001f0dd9";
		wait for Clk_period;
		Addr <=  "00001101110101";
		Trees_din <= x"00980dd9";
		wait for Clk_period;
		Addr <=  "00001101110110";
		Trees_din <= x"000ec834";
		wait for Clk_period;
		Addr <=  "00001101110111";
		Trees_din <= x"00054904";
		wait for Clk_period;
		Addr <=  "00001101111000";
		Trees_din <= x"ff7e0e55";
		wait for Clk_period;
		Addr <=  "00001101111001";
		Trees_din <= x"15fa6f14";
		wait for Clk_period;
		Addr <=  "00001101111010";
		Trees_din <= x"0b03b210";
		wait for Clk_period;
		Addr <=  "00001101111011";
		Trees_din <= x"19009208";
		wait for Clk_period;
		Addr <=  "00001101111100";
		Trees_din <= x"05072404";
		wait for Clk_period;
		Addr <=  "00001101111101";
		Trees_din <= x"00050e55";
		wait for Clk_period;
		Addr <=  "00001101111110";
		Trees_din <= x"ffac0e55";
		wait for Clk_period;
		Addr <=  "00001101111111";
		Trees_din <= x"0501ea04";
		wait for Clk_period;
		Addr <=  "00001110000000";
		Trees_din <= x"000c0e55";
		wait for Clk_period;
		Addr <=  "00001110000001";
		Trees_din <= x"00420e55";
		wait for Clk_period;
		Addr <=  "00001110000010";
		Trees_din <= x"ff5a0e55";
		wait for Clk_period;
		Addr <=  "00001110000011";
		Trees_din <= x"03fd4610";
		wait for Clk_period;
		Addr <=  "00001110000100";
		Trees_din <= x"0b00ae08";
		wait for Clk_period;
		Addr <=  "00001110000101";
		Trees_din <= x"12009804";
		wait for Clk_period;
		Addr <=  "00001110000110";
		Trees_din <= x"ff970e55";
		wait for Clk_period;
		Addr <=  "00001110000111";
		Trees_din <= x"001a0e55";
		wait for Clk_period;
		Addr <=  "00001110001000";
		Trees_din <= x"08005a04";
		wait for Clk_period;
		Addr <=  "00001110001001";
		Trees_din <= x"005c0e55";
		wait for Clk_period;
		Addr <=  "00001110001010";
		Trees_din <= x"ffc50e55";
		wait for Clk_period;
		Addr <=  "00001110001011";
		Trees_din <= x"000c1008";
		wait for Clk_period;
		Addr <=  "00001110001100";
		Trees_din <= x"09faf104";
		wait for Clk_period;
		Addr <=  "00001110001101";
		Trees_din <= x"ffe00e55";
		wait for Clk_period;
		Addr <=  "00001110001110";
		Trees_din <= x"003e0e55";
		wait for Clk_period;
		Addr <=  "00001110001111";
		Trees_din <= x"007b0e55";
		wait for Clk_period;
		Addr <=  "00001110010000";
		Trees_din <= x"09f71e04";
		wait for Clk_period;
		Addr <=  "00001110010001";
		Trees_din <= x"00180e55";
		wait for Clk_period;
		Addr <=  "00001110010010";
		Trees_din <= x"05f92504";
		wait for Clk_period;
		Addr <=  "00001110010011";
		Trees_din <= x"001d0e55";
		wait for Clk_period;
		Addr <=  "00001110010100";
		Trees_din <= x"00970e55";
		wait for Clk_period;
		Addr <=  "00001110010101";
		Trees_din <= x"000ec838";
		wait for Clk_period;
		Addr <=  "00001110010110";
		Trees_din <= x"000b0b18";
		wait for Clk_period;
		Addr <=  "00001110010111";
		Trees_din <= x"01fb660c";
		wait for Clk_period;
		Addr <=  "00001110011000";
		Trees_din <= x"07005304";
		wait for Clk_period;
		Addr <=  "00001110011001";
		Trees_din <= x"00290ed9";
		wait for Clk_period;
		Addr <=  "00001110011010";
		Trees_din <= x"0507e104";
		wait for Clk_period;
		Addr <=  "00001110011011";
		Trees_din <= x"fffe0ed9";
		wait for Clk_period;
		Addr <=  "00001110011100";
		Trees_din <= x"ffa90ed9";
		wait for Clk_period;
		Addr <=  "00001110011101";
		Trees_din <= x"07005b08";
		wait for Clk_period;
		Addr <=  "00001110011110";
		Trees_din <= x"11035704";
		wait for Clk_period;
		Addr <=  "00001110011111";
		Trees_din <= x"ff830ed9";
		wait for Clk_period;
		Addr <=  "00001110100000";
		Trees_din <= x"ffdf0ed9";
		wait for Clk_period;
		Addr <=  "00001110100001";
		Trees_din <= x"ffea0ed9";
		wait for Clk_period;
		Addr <=  "00001110100010";
		Trees_din <= x"1c003810";
		wait for Clk_period;
		Addr <=  "00001110100011";
		Trees_din <= x"0f00d90c";
		wait for Clk_period;
		Addr <=  "00001110100100";
		Trees_din <= x"09fa4504";
		wait for Clk_period;
		Addr <=  "00001110100101";
		Trees_din <= x"ffaa0ed9";
		wait for Clk_period;
		Addr <=  "00001110100110";
		Trees_din <= x"1900a904";
		wait for Clk_period;
		Addr <=  "00001110100111";
		Trees_din <= x"00510ed9";
		wait for Clk_period;
		Addr <=  "00001110101000";
		Trees_din <= x"fff10ed9";
		wait for Clk_period;
		Addr <=  "00001110101001";
		Trees_din <= x"00700ed9";
		wait for Clk_period;
		Addr <=  "00001110101010";
		Trees_din <= x"1e006d04";
		wait for Clk_period;
		Addr <=  "00001110101011";
		Trees_din <= x"ff3d0ed9";
		wait for Clk_period;
		Addr <=  "00001110101100";
		Trees_din <= x"06fc5e04";
		wait for Clk_period;
		Addr <=  "00001110101101";
		Trees_din <= x"ffcb0ed9";
		wait for Clk_period;
		Addr <=  "00001110101110";
		Trees_din <= x"03fbf704";
		wait for Clk_period;
		Addr <=  "00001110101111";
		Trees_din <= x"fff10ed9";
		wait for Clk_period;
		Addr <=  "00001110110000";
		Trees_din <= x"006e0ed9";
		wait for Clk_period;
		Addr <=  "00001110110001";
		Trees_din <= x"0508d708";
		wait for Clk_period;
		Addr <=  "00001110110010";
		Trees_din <= x"04044704";
		wait for Clk_period;
		Addr <=  "00001110110011";
		Trees_din <= x"00950ed9";
		wait for Clk_period;
		Addr <=  "00001110110100";
		Trees_din <= x"00130ed9";
		wait for Clk_period;
		Addr <=  "00001110110101";
		Trees_din <= x"00110ed9";
		wait for Clk_period;
		Addr <=  "00001110110110";
		Trees_din <= x"000ec838";
		wait for Clk_period;
		Addr <=  "00001110110111";
		Trees_din <= x"00054904";
		wait for Clk_period;
		Addr <=  "00001110111000";
		Trees_din <= x"ff870f5d";
		wait for Clk_period;
		Addr <=  "00001110111001";
		Trees_din <= x"0a013218";
		wait for Clk_period;
		Addr <=  "00001110111010";
		Trees_din <= x"000a0708";
		wait for Clk_period;
		Addr <=  "00001110111011";
		Trees_din <= x"02041304";
		wait for Clk_period;
		Addr <=  "00001110111100";
		Trees_din <= x"ffc20f5d";
		wait for Clk_period;
		Addr <=  "00001110111101";
		Trees_din <= x"00040f5d";
		wait for Clk_period;
		Addr <=  "00001110111110";
		Trees_din <= x"0c006608";
		wait for Clk_period;
		Addr <=  "00001110111111";
		Trees_din <= x"1a004d04";
		wait for Clk_period;
		Addr <=  "00001111000000";
		Trees_din <= x"ffdc0f5d";
		wait for Clk_period;
		Addr <=  "00001111000001";
		Trees_din <= x"003f0f5d";
		wait for Clk_period;
		Addr <=  "00001111000010";
		Trees_din <= x"05098d04";
		wait for Clk_period;
		Addr <=  "00001111000011";
		Trees_din <= x"00710f5d";
		wait for Clk_period;
		Addr <=  "00001111000100";
		Trees_din <= x"00270f5d";
		wait for Clk_period;
		Addr <=  "00001111000101";
		Trees_din <= x"10028710";
		wait for Clk_period;
		Addr <=  "00001111000110";
		Trees_din <= x"0a028908";
		wait for Clk_period;
		Addr <=  "00001111000111";
		Trees_din <= x"01fabf04";
		wait for Clk_period;
		Addr <=  "00001111001000";
		Trees_din <= x"00220f5d";
		wait for Clk_period;
		Addr <=  "00001111001001";
		Trees_din <= x"ffc00f5d";
		wait for Clk_period;
		Addr <=  "00001111001010";
		Trees_din <= x"01fa9d04";
		wait for Clk_period;
		Addr <=  "00001111001011";
		Trees_din <= x"000d0f5d";
		wait for Clk_period;
		Addr <=  "00001111001100";
		Trees_din <= x"004f0f5d";
		wait for Clk_period;
		Addr <=  "00001111001101";
		Trees_din <= x"08005408";
		wait for Clk_period;
		Addr <=  "00001111001110";
		Trees_din <= x"1d00da04";
		wait for Clk_period;
		Addr <=  "00001111001111";
		Trees_din <= x"ff480f5d";
		wait for Clk_period;
		Addr <=  "00001111010000";
		Trees_din <= x"ffd30f5d";
		wait for Clk_period;
		Addr <=  "00001111010001";
		Trees_din <= x"00080f5d";
		wait for Clk_period;
		Addr <=  "00001111010010";
		Trees_din <= x"0508d708";
		wait for Clk_period;
		Addr <=  "00001111010011";
		Trees_din <= x"04044704";
		wait for Clk_period;
		Addr <=  "00001111010100";
		Trees_din <= x"00940f5d";
		wait for Clk_period;
		Addr <=  "00001111010101";
		Trees_din <= x"00110f5d";
		wait for Clk_period;
		Addr <=  "00001111010110";
		Trees_din <= x"000f0f5d";
		wait for Clk_period;
		Addr <=  "00001111010111";
		Trees_din <= x"000ec838";
		wait for Clk_period;
		Addr <=  "00001111011000";
		Trees_din <= x"00087608";
		wait for Clk_period;
		Addr <=  "00001111011001";
		Trees_din <= x"11035304";
		wait for Clk_period;
		Addr <=  "00001111011010";
		Trees_din <= x"ff900fe1";
		wait for Clk_period;
		Addr <=  "00001111011011";
		Trees_din <= x"ffef0fe1";
		wait for Clk_period;
		Addr <=  "00001111011100";
		Trees_din <= x"0a013214";
		wait for Clk_period;
		Addr <=  "00001111011101";
		Trees_din <= x"0a001408";
		wait for Clk_period;
		Addr <=  "00001111011110";
		Trees_din <= x"08005104";
		wait for Clk_period;
		Addr <=  "00001111011111";
		Trees_din <= x"00290fe1";
		wait for Clk_period;
		Addr <=  "00001111100000";
		Trees_din <= x"ffcf0fe1";
		wait for Clk_period;
		Addr <=  "00001111100001";
		Trees_din <= x"0ffeb104";
		wait for Clk_period;
		Addr <=  "00001111100010";
		Trees_din <= x"fff30fe1";
		wait for Clk_period;
		Addr <=  "00001111100011";
		Trees_din <= x"13fafb04";
		wait for Clk_period;
		Addr <=  "00001111100100";
		Trees_din <= x"000d0fe1";
		wait for Clk_period;
		Addr <=  "00001111100101";
		Trees_din <= x"00700fe1";
		wait for Clk_period;
		Addr <=  "00001111100110";
		Trees_din <= x"10028710";
		wait for Clk_period;
		Addr <=  "00001111100111";
		Trees_din <= x"0d021808";
		wait for Clk_period;
		Addr <=  "00001111101000";
		Trees_din <= x"02ff9b04";
		wait for Clk_period;
		Addr <=  "00001111101001";
		Trees_din <= x"ffa80fe1";
		wait for Clk_period;
		Addr <=  "00001111101010";
		Trees_din <= x"fffe0fe1";
		wait for Clk_period;
		Addr <=  "00001111101011";
		Trees_din <= x"1e007b04";
		wait for Clk_period;
		Addr <=  "00001111101100";
		Trees_din <= x"00530fe1";
		wait for Clk_period;
		Addr <=  "00001111101101";
		Trees_din <= x"ffdb0fe1";
		wait for Clk_period;
		Addr <=  "00001111101110";
		Trees_din <= x"08005408";
		wait for Clk_period;
		Addr <=  "00001111101111";
		Trees_din <= x"1d00d904";
		wait for Clk_period;
		Addr <=  "00001111110000";
		Trees_din <= x"ff5f0fe1";
		wait for Clk_period;
		Addr <=  "00001111110001";
		Trees_din <= x"ffd80fe1";
		wait for Clk_period;
		Addr <=  "00001111110010";
		Trees_din <= x"00090fe1";
		wait for Clk_period;
		Addr <=  "00001111110011";
		Trees_din <= x"03fc0304";
		wait for Clk_period;
		Addr <=  "00001111110100";
		Trees_din <= x"001c0fe1";
		wait for Clk_period;
		Addr <=  "00001111110101";
		Trees_din <= x"0bf98b04";
		wait for Clk_period;
		Addr <=  "00001111110110";
		Trees_din <= x"00200fe1";
		wait for Clk_period;
		Addr <=  "00001111110111";
		Trees_din <= x"00920fe1";
		wait for Clk_period;
		Addr <=  "00001111111000";
		Trees_din <= x"000ec828";
		wait for Clk_period;
		Addr <=  "00001111111001";
		Trees_din <= x"00054904";
		wait for Clk_period;
		Addr <=  "00001111111010";
		Trees_din <= x"ff901045";
		wait for Clk_period;
		Addr <=  "00001111111011";
		Trees_din <= x"15fa9f0c";
		wait for Clk_period;
		Addr <=  "00001111111100";
		Trees_din <= x"16006908";
		wait for Clk_period;
		Addr <=  "00001111111101";
		Trees_din <= x"11026a04";
		wait for Clk_period;
		Addr <=  "00001111111110";
		Trees_din <= x"fff91045";
		wait for Clk_period;
		Addr <=  "00001111111111";
		Trees_din <= x"ff881045";
		wait for Clk_period;
		Addr <=  "00010000000000";
		Trees_din <= x"00181045";
		wait for Clk_period;
		Addr <=  "00010000000001";
		Trees_din <= x"1102c810";
		wait for Clk_period;
		Addr <=  "00010000000010";
		Trees_din <= x"06fe1f08";
		wait for Clk_period;
		Addr <=  "00010000000011";
		Trees_din <= x"08005304";
		wait for Clk_period;
		Addr <=  "00010000000100";
		Trees_din <= x"00441045";
		wait for Clk_period;
		Addr <=  "00010000000101";
		Trees_din <= x"fff01045";
		wait for Clk_period;
		Addr <=  "00010000000110";
		Trees_din <= x"03fd4004";
		wait for Clk_period;
		Addr <=  "00010000000111";
		Trees_din <= x"ffa51045";
		wait for Clk_period;
		Addr <=  "00010000001000";
		Trees_din <= x"00141045";
		wait for Clk_period;
		Addr <=  "00010000001001";
		Trees_din <= x"04fe2204";
		wait for Clk_period;
		Addr <=  "00010000001010";
		Trees_din <= x"00171045";
		wait for Clk_period;
		Addr <=  "00010000001011";
		Trees_din <= x"005c1045";
		wait for Clk_period;
		Addr <=  "00010000001100";
		Trees_din <= x"03fc0304";
		wait for Clk_period;
		Addr <=  "00010000001101";
		Trees_din <= x"00181045";
		wait for Clk_period;
		Addr <=  "00010000001110";
		Trees_din <= x"0bf98b04";
		wait for Clk_period;
		Addr <=  "00010000001111";
		Trees_din <= x"001c1045";
		wait for Clk_period;
		Addr <=  "00010000010000";
		Trees_din <= x"008f1045";
		wait for Clk_period;
		Addr <=  "00010000010001";
		Trees_din <= x"000ec828";
		wait for Clk_period;
		Addr <=  "00010000010010";
		Trees_din <= x"000b0b0c";
		wait for Clk_period;
		Addr <=  "00010000010011";
		Trees_din <= x"01fb6608";
		wait for Clk_period;
		Addr <=  "00010000010100";
		Trees_din <= x"0904ba04";
		wait for Clk_period;
		Addr <=  "00010000010101";
		Trees_din <= x"ffd110a9";
		wait for Clk_period;
		Addr <=  "00010000010110";
		Trees_din <= x"002a10a9";
		wait for Clk_period;
		Addr <=  "00010000010111";
		Trees_din <= x"ffa210a9";
		wait for Clk_period;
		Addr <=  "00010000011000";
		Trees_din <= x"1c00380c";
		wait for Clk_period;
		Addr <=  "00010000011001";
		Trees_din <= x"0f00d908";
		wait for Clk_period;
		Addr <=  "00010000011010";
		Trees_din <= x"0902c204";
		wait for Clk_period;
		Addr <=  "00010000011011";
		Trees_din <= x"ffc210a9";
		wait for Clk_period;
		Addr <=  "00010000011100";
		Trees_din <= x"001810a9";
		wait for Clk_period;
		Addr <=  "00010000011101";
		Trees_din <= x"006010a9";
		wait for Clk_period;
		Addr <=  "00010000011110";
		Trees_din <= x"1c003a04";
		wait for Clk_period;
		Addr <=  "00010000011111";
		Trees_din <= x"ff7810a9";
		wait for Clk_period;
		Addr <=  "00010000100000";
		Trees_din <= x"06fc5e04";
		wait for Clk_period;
		Addr <=  "00010000100001";
		Trees_din <= x"ffd210a9";
		wait for Clk_period;
		Addr <=  "00010000100010";
		Trees_din <= x"03fbf704";
		wait for Clk_period;
		Addr <=  "00010000100011";
		Trees_din <= x"fff710a9";
		wait for Clk_period;
		Addr <=  "00010000100100";
		Trees_din <= x"005a10a9";
		wait for Clk_period;
		Addr <=  "00010000100101";
		Trees_din <= x"1e008a08";
		wait for Clk_period;
		Addr <=  "00010000100110";
		Trees_din <= x"0d003504";
		wait for Clk_period;
		Addr <=  "00010000100111";
		Trees_din <= x"001f10a9";
		wait for Clk_period;
		Addr <=  "00010000101000";
		Trees_din <= x"008c10a9";
		wait for Clk_period;
		Addr <=  "00010000101001";
		Trees_din <= x"002410a9";
		wait for Clk_period;
		Addr <=  "00010000101010";
		Trees_din <= x"000ec828";
		wait for Clk_period;
		Addr <=  "00010000101011";
		Trees_din <= x"00087608";
		wait for Clk_period;
		Addr <=  "00010000101100";
		Trees_din <= x"01fc4704";
		wait for Clk_period;
		Addr <=  "00010000101101";
		Trees_din <= x"ffe7110d";
		wait for Clk_period;
		Addr <=  "00010000101110";
		Trees_din <= x"ff98110d";
		wait for Clk_period;
		Addr <=  "00010000101111";
		Trees_din <= x"03fde218";
		wait for Clk_period;
		Addr <=  "00010000110000";
		Trees_din <= x"0a01320c";
		wait for Clk_period;
		Addr <=  "00010000110001";
		Trees_din <= x"06fcfd04";
		wait for Clk_period;
		Addr <=  "00010000110010";
		Trees_din <= x"0044110d";
		wait for Clk_period;
		Addr <=  "00010000110011";
		Trees_din <= x"0f010004";
		wait for Clk_period;
		Addr <=  "00010000110100";
		Trees_din <= x"ffc9110d";
		wait for Clk_period;
		Addr <=  "00010000110101";
		Trees_din <= x"0011110d";
		wait for Clk_period;
		Addr <=  "00010000110110";
		Trees_din <= x"0d039608";
		wait for Clk_period;
		Addr <=  "00010000110111";
		Trees_din <= x"12009d04";
		wait for Clk_period;
		Addr <=  "00010000111000";
		Trees_din <= x"ff9f110d";
		wait for Clk_period;
		Addr <=  "00010000111001";
		Trees_din <= x"000a110d";
		wait for Clk_period;
		Addr <=  "00010000111010";
		Trees_din <= x"000e110d";
		wait for Clk_period;
		Addr <=  "00010000111011";
		Trees_din <= x"06fc0e04";
		wait for Clk_period;
		Addr <=  "00010000111100";
		Trees_din <= x"fff7110d";
		wait for Clk_period;
		Addr <=  "00010000111101";
		Trees_din <= x"0053110d";
		wait for Clk_period;
		Addr <=  "00010000111110";
		Trees_din <= x"1e008a08";
		wait for Clk_period;
		Addr <=  "00010000111111";
		Trees_din <= x"0d003504";
		wait for Clk_period;
		Addr <=  "00010001000000";
		Trees_din <= x"001c110d";
		wait for Clk_period;
		Addr <=  "00010001000001";
		Trees_din <= x"0089110d";
		wait for Clk_period;
		Addr <=  "00010001000010";
		Trees_din <= x"0020110d";
		wait for Clk_period;
		Addr <=  "00010001000011";
		Trees_din <= x"000ec824";
		wait for Clk_period;
		Addr <=  "00010001000100";
		Trees_din <= x"000b0b0c";
		wait for Clk_period;
		Addr <=  "00010001000101";
		Trees_din <= x"01fb6608";
		wait for Clk_period;
		Addr <=  "00010001000110";
		Trees_din <= x"0203cd04";
		wait for Clk_period;
		Addr <=  "00010001000111";
		Trees_din <= x"ffd21169";
		wait for Clk_period;
		Addr <=  "00010001001000";
		Trees_din <= x"00231169";
		wait for Clk_period;
		Addr <=  "00010001001001";
		Trees_din <= x"ffab1169";
		wait for Clk_period;
		Addr <=  "00010001001010";
		Trees_din <= x"01fcd510";
		wait for Clk_period;
		Addr <=  "00010001001011";
		Trees_din <= x"03fddd0c";
		wait for Clk_period;
		Addr <=  "00010001001100";
		Trees_din <= x"04fdec04";
		wait for Clk_period;
		Addr <=  "00010001001101";
		Trees_din <= x"00281169";
		wait for Clk_period;
		Addr <=  "00010001001110";
		Trees_din <= x"0d01c404";
		wait for Clk_period;
		Addr <=  "00010001001111";
		Trees_din <= x"00031169";
		wait for Clk_period;
		Addr <=  "00010001010000";
		Trees_din <= x"ff9a1169";
		wait for Clk_period;
		Addr <=  "00010001010001";
		Trees_din <= x"003f1169";
		wait for Clk_period;
		Addr <=  "00010001010010";
		Trees_din <= x"000c1004";
		wait for Clk_period;
		Addr <=  "00010001010011";
		Trees_din <= x"00131169";
		wait for Clk_period;
		Addr <=  "00010001010100";
		Trees_din <= x"00541169";
		wait for Clk_period;
		Addr <=  "00010001010101";
		Trees_din <= x"19007c04";
		wait for Clk_period;
		Addr <=  "00010001010110";
		Trees_din <= x"001c1169";
		wait for Clk_period;
		Addr <=  "00010001010111";
		Trees_din <= x"0a000704";
		wait for Clk_period;
		Addr <=  "00010001011000";
		Trees_din <= x"00271169";
		wait for Clk_period;
		Addr <=  "00010001011001";
		Trees_din <= x"00851169";
		wait for Clk_period;
		Addr <=  "00010001011010";
		Trees_din <= x"000fb82c";
		wait for Clk_period;
		Addr <=  "00010001011011";
		Trees_din <= x"000bb818";
		wait for Clk_period;
		Addr <=  "00010001011100";
		Trees_din <= x"01fb960c";
		wait for Clk_period;
		Addr <=  "00010001011101";
		Trees_din <= x"1504b408";
		wait for Clk_period;
		Addr <=  "00010001011110";
		Trees_din <= x"04fe6e04";
		wait for Clk_period;
		Addr <=  "00010001011111";
		Trees_din <= x"ffc011cd";
		wait for Clk_period;
		Addr <=  "00010001100000";
		Trees_din <= x"000211cd";
		wait for Clk_period;
		Addr <=  "00010001100001";
		Trees_din <= x"003a11cd";
		wait for Clk_period;
		Addr <=  "00010001100010";
		Trees_din <= x"08005504";
		wait for Clk_period;
		Addr <=  "00010001100011";
		Trees_din <= x"ffa011cd";
		wait for Clk_period;
		Addr <=  "00010001100100";
		Trees_din <= x"00097504";
		wait for Clk_period;
		Addr <=  "00010001100101";
		Trees_din <= x"ffbe11cd";
		wait for Clk_period;
		Addr <=  "00010001100110";
		Trees_din <= x"001e11cd";
		wait for Clk_period;
		Addr <=  "00010001100111";
		Trees_din <= x"02faa204";
		wait for Clk_period;
		Addr <=  "00010001101000";
		Trees_din <= x"ffc611cd";
		wait for Clk_period;
		Addr <=  "00010001101001";
		Trees_din <= x"13028708";
		wait for Clk_period;
		Addr <=  "00010001101010";
		Trees_din <= x"1d00b104";
		wait for Clk_period;
		Addr <=  "00010001101011";
		Trees_din <= x"fffa11cd";
		wait for Clk_period;
		Addr <=  "00010001101100";
		Trees_din <= x"005911cd";
		wait for Clk_period;
		Addr <=  "00010001101101";
		Trees_din <= x"10019d04";
		wait for Clk_period;
		Addr <=  "00010001101110";
		Trees_din <= x"001d11cd";
		wait for Clk_period;
		Addr <=  "00010001101111";
		Trees_din <= x"ffbc11cd";
		wait for Clk_period;
		Addr <=  "00010001110000";
		Trees_din <= x"09f99904";
		wait for Clk_period;
		Addr <=  "00010001110001";
		Trees_din <= x"001d11cd";
		wait for Clk_period;
		Addr <=  "00010001110010";
		Trees_din <= x"008211cd";
		wait for Clk_period;
		Addr <=  "00010001110011";
		Trees_din <= x"000ec82c";
		wait for Clk_period;
		Addr <=  "00010001110100";
		Trees_din <= x"0007ff08";
		wait for Clk_period;
		Addr <=  "00010001110101";
		Trees_din <= x"01fc1904";
		wait for Clk_period;
		Addr <=  "00010001110110";
		Trees_din <= x"ffea1231";
		wait for Clk_period;
		Addr <=  "00010001110111";
		Trees_din <= x"ffa51231";
		wait for Clk_period;
		Addr <=  "00010001111000";
		Trees_din <= x"03fde21c";
		wait for Clk_period;
		Addr <=  "00010001111001";
		Trees_din <= x"09fbe00c";
		wait for Clk_period;
		Addr <=  "00010001111010";
		Trees_din <= x"13fcd504";
		wait for Clk_period;
		Addr <=  "00010001111011";
		Trees_din <= x"004a1231";
		wait for Clk_period;
		Addr <=  "00010001111100";
		Trees_din <= x"0a01d104";
		wait for Clk_period;
		Addr <=  "00010001111101";
		Trees_din <= x"000f1231";
		wait for Clk_period;
		Addr <=  "00010001111110";
		Trees_din <= x"ffca1231";
		wait for Clk_period;
		Addr <=  "00010001111111";
		Trees_din <= x"10027808";
		wait for Clk_period;
		Addr <=  "00010010000000";
		Trees_din <= x"0904f604";
		wait for Clk_period;
		Addr <=  "00010010000001";
		Trees_din <= x"00231231";
		wait for Clk_period;
		Addr <=  "00010010000010";
		Trees_din <= x"ffcc1231";
		wait for Clk_period;
		Addr <=  "00010010000011";
		Trees_din <= x"0f028704";
		wait for Clk_period;
		Addr <=  "00010010000100";
		Trees_din <= x"ffe61231";
		wait for Clk_period;
		Addr <=  "00010010000101";
		Trees_din <= x"ff991231";
		wait for Clk_period;
		Addr <=  "00010010000110";
		Trees_din <= x"13fc3704";
		wait for Clk_period;
		Addr <=  "00010010000111";
		Trees_din <= x"fff01231";
		wait for Clk_period;
		Addr <=  "00010010001000";
		Trees_din <= x"004c1231";
		wait for Clk_period;
		Addr <=  "00010010001001";
		Trees_din <= x"02ff2a04";
		wait for Clk_period;
		Addr <=  "00010010001010";
		Trees_din <= x"007c1231";
		wait for Clk_period;
		Addr <=  "00010010001011";
		Trees_din <= x"002e1231";
		wait for Clk_period;
		Addr <=  "00010010001100";
		Trees_din <= x"000fb824";
		wait for Clk_period;
		Addr <=  "00010010001101";
		Trees_din <= x"000c1014";
		wait for Clk_period;
		Addr <=  "00010010001110";
		Trees_din <= x"08004b04";
		wait for Clk_period;
		Addr <=  "00010010001111";
		Trees_din <= x"0010127d";
		wait for Clk_period;
		Addr <=  "00010010010000";
		Trees_din <= x"1103530c";
		wait for Clk_period;
		Addr <=  "00010010010001";
		Trees_din <= x"0fff1104";
		wait for Clk_period;
		Addr <=  "00010010010010";
		Trees_din <= x"fff3127d";
		wait for Clk_period;
		Addr <=  "00010010010011";
		Trees_din <= x"14014004";
		wait for Clk_period;
		Addr <=  "00010010010100";
		Trees_din <= x"ffe8127d";
		wait for Clk_period;
		Addr <=  "00010010010101";
		Trees_din <= x"ffa5127d";
		wait for Clk_period;
		Addr <=  "00010010010110";
		Trees_din <= x"0002127d";
		wait for Clk_period;
		Addr <=  "00010010010111";
		Trees_din <= x"02faa204";
		wait for Clk_period;
		Addr <=  "00010010011000";
		Trees_din <= x"ffce127d";
		wait for Clk_period;
		Addr <=  "00010010011001";
		Trees_din <= x"13028708";
		wait for Clk_period;
		Addr <=  "00010010011010";
		Trees_din <= x"08005904";
		wait for Clk_period;
		Addr <=  "00010010011011";
		Trees_din <= x"0056127d";
		wait for Clk_period;
		Addr <=  "00010010011100";
		Trees_din <= x"fffe127d";
		wait for Clk_period;
		Addr <=  "00010010011101";
		Trees_din <= x"ffeb127d";
		wait for Clk_period;
		Addr <=  "00010010011110";
		Trees_din <= x"006e127d";
		wait for Clk_period;
		Addr <=  "00010010011111";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00010010100000";
		Trees_din <= x"000fb828";
		wait for Clk_period;
		Addr <=  "00010010100001";
		Trees_din <= x"000c1014";
		wait for Clk_period;
		Addr <=  "00010010100010";
		Trees_din <= x"07005408";
		wait for Clk_period;
		Addr <=  "00010010100011";
		Trees_din <= x"0c00cc04";
		wait for Clk_period;
		Addr <=  "00010010100100";
		Trees_din <= x"003312d5";
		wait for Clk_period;
		Addr <=  "00010010100101";
		Trees_din <= x"ffd412d5";
		wait for Clk_period;
		Addr <=  "00010010100110";
		Trees_din <= x"0c00c904";
		wait for Clk_period;
		Addr <=  "00010010100111";
		Trees_din <= x"ffb212d5";
		wait for Clk_period;
		Addr <=  "00010010101000";
		Trees_din <= x"07005704";
		wait for Clk_period;
		Addr <=  "00010010101001";
		Trees_din <= x"ffc712d5";
		wait for Clk_period;
		Addr <=  "00010010101010";
		Trees_din <= x"001512d5";
		wait for Clk_period;
		Addr <=  "00010010101011";
		Trees_din <= x"07005408";
		wait for Clk_period;
		Addr <=  "00010010101100";
		Trees_din <= x"02fbe804";
		wait for Clk_period;
		Addr <=  "00010010101101";
		Trees_din <= x"ffb612d5";
		wait for Clk_period;
		Addr <=  "00010010101110";
		Trees_din <= x"001512d5";
		wait for Clk_period;
		Addr <=  "00010010101111";
		Trees_din <= x"13028708";
		wait for Clk_period;
		Addr <=  "00010010110000";
		Trees_din <= x"08005904";
		wait for Clk_period;
		Addr <=  "00010010110001";
		Trees_din <= x"006212d5";
		wait for Clk_period;
		Addr <=  "00010010110010";
		Trees_din <= x"fffe12d5";
		wait for Clk_period;
		Addr <=  "00010010110011";
		Trees_din <= x"ffe912d5";
		wait for Clk_period;
		Addr <=  "00010010110100";
		Trees_din <= x"006812d5";
		wait for Clk_period;
		Addr <=  "00010010110101";
		Trees_din <= x"000ec824";
		wait for Clk_period;
		Addr <=  "00010010110110";
		Trees_din <= x"0007ff04";
		wait for Clk_period;
		Addr <=  "00010010110111";
		Trees_din <= x"ffb91329";
		wait for Clk_period;
		Addr <=  "00010010111000";
		Trees_din <= x"15fa9f08";
		wait for Clk_period;
		Addr <=  "00010010111001";
		Trees_din <= x"11026a04";
		wait for Clk_period;
		Addr <=  "00010010111010";
		Trees_din <= x"000b1329";
		wait for Clk_period;
		Addr <=  "00010010111011";
		Trees_din <= x"ffb61329";
		wait for Clk_period;
		Addr <=  "00010010111100";
		Trees_din <= x"03fd4610";
		wait for Clk_period;
		Addr <=  "00010010111101";
		Trees_din <= x"0b004208";
		wait for Clk_period;
		Addr <=  "00010010111110";
		Trees_din <= x"18003604";
		wait for Clk_period;
		Addr <=  "00010010111111";
		Trees_din <= x"ffff1329";
		wait for Clk_period;
		Addr <=  "00010011000000";
		Trees_din <= x"ffc01329";
		wait for Clk_period;
		Addr <=  "00010011000001";
		Trees_din <= x"13fcd504";
		wait for Clk_period;
		Addr <=  "00010011000010";
		Trees_din <= x"00491329";
		wait for Clk_period;
		Addr <=  "00010011000011";
		Trees_din <= x"fff31329";
		wait for Clk_period;
		Addr <=  "00010011000100";
		Trees_din <= x"09faf104";
		wait for Clk_period;
		Addr <=  "00010011000101";
		Trees_din <= x"00041329";
		wait for Clk_period;
		Addr <=  "00010011000110";
		Trees_din <= x"00491329";
		wait for Clk_period;
		Addr <=  "00010011000111";
		Trees_din <= x"07005a04";
		wait for Clk_period;
		Addr <=  "00010011001000";
		Trees_din <= x"006e1329";
		wait for Clk_period;
		Addr <=  "00010011001001";
		Trees_din <= x"00191329";
		wait for Clk_period;
		Addr <=  "00010011001010";
		Trees_din <= x"000c1010";
		wait for Clk_period;
		Addr <=  "00010011001011";
		Trees_din <= x"01fb9608";
		wait for Clk_period;
		Addr <=  "00010011001100";
		Trees_din <= x"1000ae04";
		wait for Clk_period;
		Addr <=  "00010011001101";
		Trees_din <= x"00231375";
		wait for Clk_period;
		Addr <=  "00010011001110";
		Trees_din <= x"ffd81375";
		wait for Clk_period;
		Addr <=  "00010011001111";
		Trees_din <= x"08005504";
		wait for Clk_period;
		Addr <=  "00010011010000";
		Trees_din <= x"ffaf1375";
		wait for Clk_period;
		Addr <=  "00010011010001";
		Trees_din <= x"fff41375";
		wait for Clk_period;
		Addr <=  "00010011010010";
		Trees_din <= x"03fdea14";
		wait for Clk_period;
		Addr <=  "00010011010011";
		Trees_din <= x"0d01fb08";
		wait for Clk_period;
		Addr <=  "00010011010100";
		Trees_din <= x"06fdb404";
		wait for Clk_period;
		Addr <=  "00010011010101";
		Trees_din <= x"004b1375";
		wait for Clk_period;
		Addr <=  "00010011010110";
		Trees_din <= x"fffd1375";
		wait for Clk_period;
		Addr <=  "00010011010111";
		Trees_din <= x"0d034b08";
		wait for Clk_period;
		Addr <=  "00010011011000";
		Trees_din <= x"19008f04";
		wait for Clk_period;
		Addr <=  "00010011011001";
		Trees_din <= x"ffb11375";
		wait for Clk_period;
		Addr <=  "00010011011010";
		Trees_din <= x"fff51375";
		wait for Clk_period;
		Addr <=  "00010011011011";
		Trees_din <= x"00261375";
		wait for Clk_period;
		Addr <=  "00010011011100";
		Trees_din <= x"006a1375";
		wait for Clk_period;
		Addr <=  "00010011011101";
		Trees_din <= x"000fb824";
		wait for Clk_period;
		Addr <=  "00010011011110";
		Trees_din <= x"000a0708";
		wait for Clk_period;
		Addr <=  "00010011011111";
		Trees_din <= x"01fb6604";
		wait for Clk_period;
		Addr <=  "00010011100000";
		Trees_din <= x"fff213c1";
		wait for Clk_period;
		Addr <=  "00010011100001";
		Trees_din <= x"ffb513c1";
		wait for Clk_period;
		Addr <=  "00010011100010";
		Trees_din <= x"0a013b0c";
		wait for Clk_period;
		Addr <=  "00010011100011";
		Trees_din <= x"0a001404";
		wait for Clk_period;
		Addr <=  "00010011100100";
		Trees_din <= x"ffed13c1";
		wait for Clk_period;
		Addr <=  "00010011100101";
		Trees_din <= x"01fabf04";
		wait for Clk_period;
		Addr <=  "00010011100110";
		Trees_din <= x"000413c1";
		wait for Clk_period;
		Addr <=  "00010011100111";
		Trees_din <= x"005a13c1";
		wait for Clk_period;
		Addr <=  "00010011101000";
		Trees_din <= x"08005308";
		wait for Clk_period;
		Addr <=  "00010011101001";
		Trees_din <= x"1c003804";
		wait for Clk_period;
		Addr <=  "00010011101010";
		Trees_din <= x"fffb13c1";
		wait for Clk_period;
		Addr <=  "00010011101011";
		Trees_din <= x"ffab13c1";
		wait for Clk_period;
		Addr <=  "00010011101100";
		Trees_din <= x"05079604";
		wait for Clk_period;
		Addr <=  "00010011101101";
		Trees_din <= x"003e13c1";
		wait for Clk_period;
		Addr <=  "00010011101110";
		Trees_din <= x"ffdf13c1";
		wait for Clk_period;
		Addr <=  "00010011101111";
		Trees_din <= x"005913c1";
		wait for Clk_period;
		Addr <=  "00010011110000";
		Trees_din <= x"000c1014";
		wait for Clk_period;
		Addr <=  "00010011110001";
		Trees_din <= x"07005408";
		wait for Clk_period;
		Addr <=  "00010011110010";
		Trees_din <= x"01fb9604";
		wait for Clk_period;
		Addr <=  "00010011110011";
		Trees_din <= x"00211415";
		wait for Clk_period;
		Addr <=  "00010011110100";
		Trees_din <= x"ffda1415";
		wait for Clk_period;
		Addr <=  "00010011110101";
		Trees_din <= x"0c00c904";
		wait for Clk_period;
		Addr <=  "00010011110110";
		Trees_din <= x"ffb91415";
		wait for Clk_period;
		Addr <=  "00010011110111";
		Trees_din <= x"0a00e004";
		wait for Clk_period;
		Addr <=  "00010011111000";
		Trees_din <= x"000e1415";
		wait for Clk_period;
		Addr <=  "00010011111001";
		Trees_din <= x"ffd81415";
		wait for Clk_period;
		Addr <=  "00010011111010";
		Trees_din <= x"03fdea14";
		wait for Clk_period;
		Addr <=  "00010011111011";
		Trees_din <= x"0d01fb08";
		wait for Clk_period;
		Addr <=  "00010011111100";
		Trees_din <= x"06fdb404";
		wait for Clk_period;
		Addr <=  "00010011111101";
		Trees_din <= x"00451415";
		wait for Clk_period;
		Addr <=  "00010011111110";
		Trees_din <= x"fffa1415";
		wait for Clk_period;
		Addr <=  "00010011111111";
		Trees_din <= x"0d034b08";
		wait for Clk_period;
		Addr <=  "00010100000000";
		Trees_din <= x"19008f04";
		wait for Clk_period;
		Addr <=  "00010100000001";
		Trees_din <= x"ffb91415";
		wait for Clk_period;
		Addr <=  "00010100000010";
		Trees_din <= x"fff61415";
		wait for Clk_period;
		Addr <=  "00010100000011";
		Trees_din <= x"00261415";
		wait for Clk_period;
		Addr <=  "00010100000100";
		Trees_din <= x"00601415";
		wait for Clk_period;
		Addr <=  "00010100000101";
		Trees_din <= x"000fb820";
		wait for Clk_period;
		Addr <=  "00010100000110";
		Trees_din <= x"000b0b0c";
		wait for Clk_period;
		Addr <=  "00010100000111";
		Trees_din <= x"07005404";
		wait for Clk_period;
		Addr <=  "00010100001000";
		Trees_din <= x"ffff1459";
		wait for Clk_period;
		Addr <=  "00010100001001";
		Trees_din <= x"07005804";
		wait for Clk_period;
		Addr <=  "00010100001010";
		Trees_din <= x"ffb41459";
		wait for Clk_period;
		Addr <=  "00010100001011";
		Trees_din <= x"fff11459";
		wait for Clk_period;
		Addr <=  "00010100001100";
		Trees_din <= x"01fcd510";
		wait for Clk_period;
		Addr <=  "00010100001101";
		Trees_din <= x"03fddd0c";
		wait for Clk_period;
		Addr <=  "00010100001110";
		Trees_din <= x"04fdec04";
		wait for Clk_period;
		Addr <=  "00010100001111";
		Trees_din <= x"00221459";
		wait for Clk_period;
		Addr <=  "00010100010000";
		Trees_din <= x"0d01dd04";
		wait for Clk_period;
		Addr <=  "00010100010001";
		Trees_din <= x"fff91459";
		wait for Clk_period;
		Addr <=  "00010100010010";
		Trees_din <= x"ffba1459";
		wait for Clk_period;
		Addr <=  "00010100010011";
		Trees_din <= x"002c1459";
		wait for Clk_period;
		Addr <=  "00010100010100";
		Trees_din <= x"002b1459";
		wait for Clk_period;
		Addr <=  "00010100010101";
		Trees_din <= x"00501459";
		wait for Clk_period;
		Addr <=  "00010100010110";
		Trees_din <= x"000e0620";
		wait for Clk_period;
		Addr <=  "00010100010111";
		Trees_din <= x"15faaf08";
		wait for Clk_period;
		Addr <=  "00010100011000";
		Trees_din <= x"0c00c704";
		wait for Clk_period;
		Addr <=  "00010100011001";
		Trees_din <= x"ffb814a5";
		wait for Clk_period;
		Addr <=  "00010100011010";
		Trees_din <= x"fff014a5";
		wait for Clk_period;
		Addr <=  "00010100011011";
		Trees_din <= x"06fcfd0c";
		wait for Clk_period;
		Addr <=  "00010100011100";
		Trees_din <= x"1504dc08";
		wait for Clk_period;
		Addr <=  "00010100011101";
		Trees_din <= x"0a012604";
		wait for Clk_period;
		Addr <=  "00010100011110";
		Trees_din <= x"004114a5";
		wait for Clk_period;
		Addr <=  "00010100011111";
		Trees_din <= x"000414a5";
		wait for Clk_period;
		Addr <=  "00010100100000";
		Trees_din <= x"ffef14a5";
		wait for Clk_period;
		Addr <=  "00010100100001";
		Trees_din <= x"1d00db08";
		wait for Clk_period;
		Addr <=  "00010100100010";
		Trees_din <= x"02026404";
		wait for Clk_period;
		Addr <=  "00010100100011";
		Trees_din <= x"002b14a5";
		wait for Clk_period;
		Addr <=  "00010100100100";
		Trees_din <= x"ffd414a5";
		wait for Clk_period;
		Addr <=  "00010100100101";
		Trees_din <= x"ffc114a5";
		wait for Clk_period;
		Addr <=  "00010100100110";
		Trees_din <= x"03fc8804";
		wait for Clk_period;
		Addr <=  "00010100100111";
		Trees_din <= x"ffef14a5";
		wait for Clk_period;
		Addr <=  "00010100101000";
		Trees_din <= x"005a14a5";
		wait for Clk_period;
		Addr <=  "00010100101001";
		Trees_din <= x"000c1010";
		wait for Clk_period;
		Addr <=  "00010100101010";
		Trees_din <= x"1505420c";
		wait for Clk_period;
		Addr <=  "00010100101011";
		Trees_din <= x"1102f908";
		wait for Clk_period;
		Addr <=  "00010100101100";
		Trees_din <= x"08005104";
		wait for Clk_period;
		Addr <=  "00010100101101";
		Trees_din <= x"fffa14e1";
		wait for Clk_period;
		Addr <=  "00010100101110";
		Trees_din <= x"ffbc14e1";
		wait for Clk_period;
		Addr <=  "00010100101111";
		Trees_din <= x"fffe14e1";
		wait for Clk_period;
		Addr <=  "00010100110000";
		Trees_din <= x"000914e1";
		wait for Clk_period;
		Addr <=  "00010100110001";
		Trees_din <= x"03fdea0c";
		wait for Clk_period;
		Addr <=  "00010100110010";
		Trees_din <= x"12009808";
		wait for Clk_period;
		Addr <=  "00010100110011";
		Trees_din <= x"1e006d04";
		wait for Clk_period;
		Addr <=  "00010100110100";
		Trees_din <= x"ffc914e1";
		wait for Clk_period;
		Addr <=  "00010100110101";
		Trees_din <= x"001914e1";
		wait for Clk_period;
		Addr <=  "00010100110110";
		Trees_din <= x"002e14e1";
		wait for Clk_period;
		Addr <=  "00010100110111";
		Trees_din <= x"005114e1";
		wait for Clk_period;
		Addr <=  "00010100111000";
		Trees_din <= x"000c1010";
		wait for Clk_period;
		Addr <=  "00010100111001";
		Trees_din <= x"01fb9608";
		wait for Clk_period;
		Addr <=  "00010100111010";
		Trees_din <= x"08005204";
		wait for Clk_period;
		Addr <=  "00010100111011";
		Trees_din <= x"00201525";
		wait for Clk_period;
		Addr <=  "00010100111100";
		Trees_din <= x"ffdd1525";
		wait for Clk_period;
		Addr <=  "00010100111101";
		Trees_din <= x"08005504";
		wait for Clk_period;
		Addr <=  "00010100111110";
		Trees_din <= x"ffbd1525";
		wait for Clk_period;
		Addr <=  "00010100111111";
		Trees_din <= x"fff81525";
		wait for Clk_period;
		Addr <=  "00010101000000";
		Trees_din <= x"01fbc70c";
		wait for Clk_period;
		Addr <=  "00010101000001";
		Trees_din <= x"03fcf108";
		wait for Clk_period;
		Addr <=  "00010101000010";
		Trees_din <= x"0d028504";
		wait for Clk_period;
		Addr <=  "00010101000011";
		Trees_din <= x"00011525";
		wait for Clk_period;
		Addr <=  "00010101000100";
		Trees_din <= x"ffcd1525";
		wait for Clk_period;
		Addr <=  "00010101000101";
		Trees_din <= x"00271525";
		wait for Clk_period;
		Addr <=  "00010101000110";
		Trees_din <= x"08005604";
		wait for Clk_period;
		Addr <=  "00010101000111";
		Trees_din <= x"00531525";
		wait for Clk_period;
		Addr <=  "00010101001000";
		Trees_din <= x"00181525";
		wait for Clk_period;
		Addr <=  "00010101001001";
		Trees_din <= x"000e0618";
		wait for Clk_period;
		Addr <=  "00010101001010";
		Trees_din <= x"15faaf04";
		wait for Clk_period;
		Addr <=  "00010101001011";
		Trees_din <= x"ffca1561";
		wait for Clk_period;
		Addr <=  "00010101001100";
		Trees_din <= x"06fcfd08";
		wait for Clk_period;
		Addr <=  "00010101001101";
		Trees_din <= x"1503c304";
		wait for Clk_period;
		Addr <=  "00010101001110";
		Trees_din <= x"00381561";
		wait for Clk_period;
		Addr <=  "00010101001111";
		Trees_din <= x"fffb1561";
		wait for Clk_period;
		Addr <=  "00010101010000";
		Trees_din <= x"1d00db08";
		wait for Clk_period;
		Addr <=  "00010101010001";
		Trees_din <= x"02026404";
		wait for Clk_period;
		Addr <=  "00010101010010";
		Trees_din <= x"00271561";
		wait for Clk_period;
		Addr <=  "00010101010011";
		Trees_din <= x"ffd81561";
		wait for Clk_period;
		Addr <=  "00010101010100";
		Trees_din <= x"ffc51561";
		wait for Clk_period;
		Addr <=  "00010101010101";
		Trees_din <= x"03fc8804";
		wait for Clk_period;
		Addr <=  "00010101010110";
		Trees_din <= x"fff51561";
		wait for Clk_period;
		Addr <=  "00010101010111";
		Trees_din <= x"004e1561";
		wait for Clk_period;
		Addr <=  "00010101011000";
		Trees_din <= x"000c100c";
		wait for Clk_period;
		Addr <=  "00010101011001";
		Trees_din <= x"07005404";
		wait for Clk_period;
		Addr <=  "00010101011010";
		Trees_din <= x"00001595";
		wait for Clk_period;
		Addr <=  "00010101011011";
		Trees_din <= x"0c00c904";
		wait for Clk_period;
		Addr <=  "00010101011100";
		Trees_din <= x"ffc21595";
		wait for Clk_period;
		Addr <=  "00010101011101";
		Trees_din <= x"fff81595";
		wait for Clk_period;
		Addr <=  "00010101011110";
		Trees_din <= x"01fbc708";
		wait for Clk_period;
		Addr <=  "00010101011111";
		Trees_din <= x"03fcf104";
		wait for Clk_period;
		Addr <=  "00010101100000";
		Trees_din <= x"ffe41595";
		wait for Clk_period;
		Addr <=  "00010101100001";
		Trees_din <= x"00221595";
		wait for Clk_period;
		Addr <=  "00010101100010";
		Trees_din <= x"19009904";
		wait for Clk_period;
		Addr <=  "00010101100011";
		Trees_din <= x"004d1595";
		wait for Clk_period;
		Addr <=  "00010101100100";
		Trees_din <= x"00121595";
		wait for Clk_period;
		Addr <=  "00010101100101";
		Trees_din <= x"000c100c";
		wait for Clk_period;
		Addr <=  "00010101100110";
		Trees_din <= x"0007ff04";
		wait for Clk_period;
		Addr <=  "00010101100111";
		Trees_din <= x"ffc815c9";
		wait for Clk_period;
		Addr <=  "00010101101000";
		Trees_din <= x"04fee804";
		wait for Clk_period;
		Addr <=  "00010101101001";
		Trees_din <= x"ffdf15c9";
		wait for Clk_period;
		Addr <=  "00010101101010";
		Trees_din <= x"001215c9";
		wait for Clk_period;
		Addr <=  "00010101101011";
		Trees_din <= x"03fdea0c";
		wait for Clk_period;
		Addr <=  "00010101101100";
		Trees_din <= x"12009808";
		wait for Clk_period;
		Addr <=  "00010101101101";
		Trees_din <= x"1e006d04";
		wait for Clk_period;
		Addr <=  "00010101101110";
		Trees_din <= x"ffce15c9";
		wait for Clk_period;
		Addr <=  "00010101101111";
		Trees_din <= x"001715c9";
		wait for Clk_period;
		Addr <=  "00010101110000";
		Trees_din <= x"002a15c9";
		wait for Clk_period;
		Addr <=  "00010101110001";
		Trees_din <= x"004515c9";
		wait for Clk_period;
		Addr <=  "00010101110010";
		Trees_din <= x"000b0b08";
		wait for Clk_period;
		Addr <=  "00010101110011";
		Trees_din <= x"0efdb104";
		wait for Clk_period;
		Addr <=  "00010101110100";
		Trees_din <= x"fffe1605";
		wait for Clk_period;
		Addr <=  "00010101110101";
		Trees_din <= x"ffcd1605";
		wait for Clk_period;
		Addr <=  "00010101110110";
		Trees_din <= x"03fdea14";
		wait for Clk_period;
		Addr <=  "00010101110111";
		Trees_din <= x"01fcd510";
		wait for Clk_period;
		Addr <=  "00010101111000";
		Trees_din <= x"01fa0c04";
		wait for Clk_period;
		Addr <=  "00010101111001";
		Trees_din <= x"00241605";
		wait for Clk_period;
		Addr <=  "00010101111010";
		Trees_din <= x"12009808";
		wait for Clk_period;
		Addr <=  "00010101111011";
		Trees_din <= x"1e006d04";
		wait for Clk_period;
		Addr <=  "00010101111100";
		Trees_din <= x"ffb41605";
		wait for Clk_period;
		Addr <=  "00010101111101";
		Trees_din <= x"fff21605";
		wait for Clk_period;
		Addr <=  "00010101111110";
		Trees_din <= x"00071605";
		wait for Clk_period;
		Addr <=  "00010101111111";
		Trees_din <= x"00251605";
		wait for Clk_period;
		Addr <=  "00010110000000";
		Trees_din <= x"00411605";
		wait for Clk_period;
		Addr <=  "00010110000001";
		Trees_din <= x"000c1010";
		wait for Clk_period;
		Addr <=  "00010110000010";
		Trees_din <= x"0fff0604";
		wait for Clk_period;
		Addr <=  "00010110000011";
		Trees_din <= x"00081639";
		wait for Clk_period;
		Addr <=  "00010110000100";
		Trees_din <= x"14014004";
		wait for Clk_period;
		Addr <=  "00010110000101";
		Trees_din <= x"fffd1639";
		wait for Clk_period;
		Addr <=  "00010110000110";
		Trees_din <= x"0d010d04";
		wait for Clk_period;
		Addr <=  "00010110000111";
		Trees_din <= x"fff41639";
		wait for Clk_period;
		Addr <=  "00010110001000";
		Trees_din <= x"ffc01639";
		wait for Clk_period;
		Addr <=  "00010110001001";
		Trees_din <= x"01fbe308";
		wait for Clk_period;
		Addr <=  "00010110001010";
		Trees_din <= x"19008f04";
		wait for Clk_period;
		Addr <=  "00010110001011";
		Trees_din <= x"ffe31639";
		wait for Clk_period;
		Addr <=  "00010110001100";
		Trees_din <= x"001e1639";
		wait for Clk_period;
		Addr <=  "00010110001101";
		Trees_din <= x"003a1639";
		wait for Clk_period;
		Addr <=  "00010110001110";
		Trees_din <= x"000fb818";
		wait for Clk_period;
		Addr <=  "00010110001111";
		Trees_din <= x"10011b0c";
		wait for Clk_period;
		Addr <=  "00010110010000";
		Trees_din <= x"16001504";
		wait for Clk_period;
		Addr <=  "00010110010001";
		Trees_din <= x"0028166d";
		wait for Clk_period;
		Addr <=  "00010110010010";
		Trees_din <= x"0a00e004";
		wait for Clk_period;
		Addr <=  "00010110010011";
		Trees_din <= x"000c166d";
		wait for Clk_period;
		Addr <=  "00010110010100";
		Trees_din <= x"ffe3166d";
		wait for Clk_period;
		Addr <=  "00010110010101";
		Trees_din <= x"1e006404";
		wait for Clk_period;
		Addr <=  "00010110010110";
		Trees_din <= x"000a166d";
		wait for Clk_period;
		Addr <=  "00010110010111";
		Trees_din <= x"09fb9604";
		wait for Clk_period;
		Addr <=  "00010110011000";
		Trees_din <= x"0005166d";
		wait for Clk_period;
		Addr <=  "00010110011001";
		Trees_din <= x"ffbc166d";
		wait for Clk_period;
		Addr <=  "00010110011010";
		Trees_din <= x"0037166d";
		wait for Clk_period;
		Addr <=  "00010110011011";
		Trees_din <= x"000c100c";
		wait for Clk_period;
		Addr <=  "00010110011100";
		Trees_din <= x"0007ff04";
		wait for Clk_period;
		Addr <=  "00010110011101";
		Trees_din <= x"ffcd16a1";
		wait for Clk_period;
		Addr <=  "00010110011110";
		Trees_din <= x"04fee804";
		wait for Clk_period;
		Addr <=  "00010110011111";
		Trees_din <= x"ffe216a1";
		wait for Clk_period;
		Addr <=  "00010110100000";
		Trees_din <= x"001016a1";
		wait for Clk_period;
		Addr <=  "00010110100001";
		Trees_din <= x"07005404";
		wait for Clk_period;
		Addr <=  "00010110100010";
		Trees_din <= x"fff416a1";
		wait for Clk_period;
		Addr <=  "00010110100011";
		Trees_din <= x"13028708";
		wait for Clk_period;
		Addr <=  "00010110100100";
		Trees_din <= x"01faa804";
		wait for Clk_period;
		Addr <=  "00010110100101";
		Trees_din <= x"000a16a1";
		wait for Clk_period;
		Addr <=  "00010110100110";
		Trees_din <= x"004916a1";
		wait for Clk_period;
		Addr <=  "00010110100111";
		Trees_din <= x"fffc16a1";
		wait for Clk_period;
		Addr <=  "00010110101000";
		Trees_din <= x"000c1010";
		wait for Clk_period;
		Addr <=  "00010110101001";
		Trees_din <= x"01fb9608";
		wait for Clk_period;
		Addr <=  "00010110101010";
		Trees_din <= x"07005404";
		wait for Clk_period;
		Addr <=  "00010110101011";
		Trees_din <= x"001c16d5";
		wait for Clk_period;
		Addr <=  "00010110101100";
		Trees_din <= x"ffe716d5";
		wait for Clk_period;
		Addr <=  "00010110101101";
		Trees_din <= x"08005504";
		wait for Clk_period;
		Addr <=  "00010110101110";
		Trees_din <= x"ffc716d5";
		wait for Clk_period;
		Addr <=  "00010110101111";
		Trees_din <= x"fffc16d5";
		wait for Clk_period;
		Addr <=  "00010110110000";
		Trees_din <= x"01fbe308";
		wait for Clk_period;
		Addr <=  "00010110110001";
		Trees_din <= x"03fcf104";
		wait for Clk_period;
		Addr <=  "00010110110010";
		Trees_din <= x"ffe916d5";
		wait for Clk_period;
		Addr <=  "00010110110011";
		Trees_din <= x"002116d5";
		wait for Clk_period;
		Addr <=  "00010110110100";
		Trees_din <= x"003316d5";
		wait for Clk_period;
		Addr <=  "00010110110101";
		Trees_din <= x"000a0704";
		wait for Clk_period;
		Addr <=  "00010110110110";
		Trees_din <= x"ffd81701";
		wait for Clk_period;
		Addr <=  "00010110110111";
		Trees_din <= x"03fdea10";
		wait for Clk_period;
		Addr <=  "00010110111000";
		Trees_din <= x"13fcf308";
		wait for Clk_period;
		Addr <=  "00010110111001";
		Trees_din <= x"06fce904";
		wait for Clk_period;
		Addr <=  "00010110111010";
		Trees_din <= x"fffb1701";
		wait for Clk_period;
		Addr <=  "00010110111011";
		Trees_din <= x"002e1701";
		wait for Clk_period;
		Addr <=  "00010110111100";
		Trees_din <= x"06fdb404";
		wait for Clk_period;
		Addr <=  "00010110111101";
		Trees_din <= x"000b1701";
		wait for Clk_period;
		Addr <=  "00010110111110";
		Trees_din <= x"ffd71701";
		wait for Clk_period;
		Addr <=  "00010110111111";
		Trees_din <= x"00341701";
		wait for Clk_period;
		Addr <=  "00010111000000";
		Trees_din <= x"000c100c";
		wait for Clk_period;
		Addr <=  "00010111000001";
		Trees_din <= x"01fb9604";
		wait for Clk_period;
		Addr <=  "00010111000010";
		Trees_din <= x"00021735";
		wait for Clk_period;
		Addr <=  "00010111000011";
		Trees_din <= x"08005504";
		wait for Clk_period;
		Addr <=  "00010111000100";
		Trees_din <= x"ffcb1735";
		wait for Clk_period;
		Addr <=  "00010111000101";
		Trees_din <= x"fffe1735";
		wait for Clk_period;
		Addr <=  "00010111000110";
		Trees_din <= x"07005404";
		wait for Clk_period;
		Addr <=  "00010111000111";
		Trees_din <= x"fff31735";
		wait for Clk_period;
		Addr <=  "00010111001000";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00010111001001";
		Trees_din <= x"003d1735";
		wait for Clk_period;
		Addr <=  "00010111001010";
		Trees_din <= x"000e6e04";
		wait for Clk_period;
		Addr <=  "00010111001011";
		Trees_din <= x"00171735";
		wait for Clk_period;
		Addr <=  "00010111001100";
		Trees_din <= x"fff61735";
		wait for Clk_period;
		Addr <=  "00010111001101";
		Trees_din <= x"000a0704";
		wait for Clk_period;
		Addr <=  "00010111001110";
		Trees_din <= x"ffda1769";
		wait for Clk_period;
		Addr <=  "00010111001111";
		Trees_din <= x"03fdea14";
		wait for Clk_period;
		Addr <=  "00010111010000";
		Trees_din <= x"0a013b08";
		wait for Clk_period;
		Addr <=  "00010111010001";
		Trees_din <= x"06fdb404";
		wait for Clk_period;
		Addr <=  "00010111010010";
		Trees_din <= x"00331769";
		wait for Clk_period;
		Addr <=  "00010111010011";
		Trees_din <= x"fff11769";
		wait for Clk_period;
		Addr <=  "00010111010100";
		Trees_din <= x"0d035708";
		wait for Clk_period;
		Addr <=  "00010111010101";
		Trees_din <= x"02ffab04";
		wait for Clk_period;
		Addr <=  "00010111010110";
		Trees_din <= x"ffc31769";
		wait for Clk_period;
		Addr <=  "00010111010111";
		Trees_din <= x"00051769";
		wait for Clk_period;
		Addr <=  "00010111011000";
		Trees_din <= x"00141769";
		wait for Clk_period;
		Addr <=  "00010111011001";
		Trees_din <= x"00301769";
		wait for Clk_period;
		Addr <=  "00010111011010";
		Trees_din <= x"000c1010";
		wait for Clk_period;
		Addr <=  "00010111011011";
		Trees_din <= x"10010f08";
		wait for Clk_period;
		Addr <=  "00010111011100";
		Trees_din <= x"01fc1904";
		wait for Clk_period;
		Addr <=  "00010111011101";
		Trees_din <= x"0012179d";
		wait for Clk_period;
		Addr <=  "00010111011110";
		Trees_din <= x"fff0179d";
		wait for Clk_period;
		Addr <=  "00010111011111";
		Trees_din <= x"08005404";
		wait for Clk_period;
		Addr <=  "00010111100000";
		Trees_din <= x"ffd0179d";
		wait for Clk_period;
		Addr <=  "00010111100001";
		Trees_din <= x"fff8179d";
		wait for Clk_period;
		Addr <=  "00010111100010";
		Trees_din <= x"15fa5e04";
		wait for Clk_period;
		Addr <=  "00010111100011";
		Trees_din <= x"fff1179d";
		wait for Clk_period;
		Addr <=  "00010111100100";
		Trees_din <= x"1301f104";
		wait for Clk_period;
		Addr <=  "00010111100101";
		Trees_din <= x"003a179d";
		wait for Clk_period;
		Addr <=  "00010111100110";
		Trees_din <= x"0007179d";
		wait for Clk_period;
		Addr <=  "00010111100111";
		Trees_din <= x"0007ff04";
		wait for Clk_period;
		Addr <=  "00010111101000";
		Trees_din <= x"ffd517d1";
		wait for Clk_period;
		Addr <=  "00010111101001";
		Trees_din <= x"03fe7c14";
		wait for Clk_period;
		Addr <=  "00010111101010";
		Trees_din <= x"12009d10";
		wait for Clk_period;
		Addr <=  "00010111101011";
		Trees_din <= x"18003a08";
		wait for Clk_period;
		Addr <=  "00010111101100";
		Trees_din <= x"03fd3604";
		wait for Clk_period;
		Addr <=  "00010111101101";
		Trees_din <= x"000117d1";
		wait for Clk_period;
		Addr <=  "00010111101110";
		Trees_din <= x"ffc117d1";
		wait for Clk_period;
		Addr <=  "00010111101111";
		Trees_din <= x"1c003f04";
		wait for Clk_period;
		Addr <=  "00010111110000";
		Trees_din <= x"003217d1";
		wait for Clk_period;
		Addr <=  "00010111110001";
		Trees_din <= x"ffe717d1";
		wait for Clk_period;
		Addr <=  "00010111110010";
		Trees_din <= x"001d17d1";
		wait for Clk_period;
		Addr <=  "00010111110011";
		Trees_din <= x"002f17d1";
		wait for Clk_period;
		Addr <=  "00010111110100";
		Trees_din <= x"000c100c";
		wait for Clk_period;
		Addr <=  "00010111110101";
		Trees_din <= x"11031e08";
		wait for Clk_period;
		Addr <=  "00010111110110";
		Trees_din <= x"06fe1a04";
		wait for Clk_period;
		Addr <=  "00010111110111";
		Trees_din <= x"fffc17fd";
		wait for Clk_period;
		Addr <=  "00010111111000";
		Trees_din <= x"ffcc17fd";
		wait for Clk_period;
		Addr <=  "00010111111001";
		Trees_din <= x"000717fd";
		wait for Clk_period;
		Addr <=  "00010111111010";
		Trees_din <= x"16000204";
		wait for Clk_period;
		Addr <=  "00010111111011";
		Trees_din <= x"fff917fd";
		wait for Clk_period;
		Addr <=  "00010111111100";
		Trees_din <= x"0b003904";
		wait for Clk_period;
		Addr <=  "00010111111101";
		Trees_din <= x"000017fd";
		wait for Clk_period;
		Addr <=  "00010111111110";
		Trees_din <= x"003917fd";
		wait for Clk_period;
		Addr <=  "00010111111111";
		Trees_din <= x"000c100c";
		wait for Clk_period;
		Addr <=  "00011000000000";
		Trees_din <= x"14014c04";
		wait for Clk_period;
		Addr <=  "00011000000001";
		Trees_din <= x"00041829";
		wait for Clk_period;
		Addr <=  "00011000000010";
		Trees_din <= x"1000e204";
		wait for Clk_period;
		Addr <=  "00011000000011";
		Trees_din <= x"fffc1829";
		wait for Clk_period;
		Addr <=  "00011000000100";
		Trees_din <= x"ffd71829";
		wait for Clk_period;
		Addr <=  "00011000000101";
		Trees_din <= x"07005404";
		wait for Clk_period;
		Addr <=  "00011000000110";
		Trees_din <= x"fff51829";
		wait for Clk_period;
		Addr <=  "00011000000111";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00011000001000";
		Trees_din <= x"00361829";
		wait for Clk_period;
		Addr <=  "00011000001001";
		Trees_din <= x"00081829";
		wait for Clk_period;
		Addr <=  "00011000001010";
		Trees_din <= x"000b0b08";
		wait for Clk_period;
		Addr <=  "00011000001011";
		Trees_din <= x"01fb6604";
		wait for Clk_period;
		Addr <=  "00011000001100";
		Trees_din <= x"00011855";
		wait for Clk_period;
		Addr <=  "00011000001101";
		Trees_din <= x"ffd71855";
		wait for Clk_period;
		Addr <=  "00011000001110";
		Trees_din <= x"1c003608";
		wait for Clk_period;
		Addr <=  "00011000001111";
		Trees_din <= x"0f00d904";
		wait for Clk_period;
		Addr <=  "00011000010000";
		Trees_din <= x"fff81855";
		wait for Clk_period;
		Addr <=  "00011000010001";
		Trees_din <= x"00481855";
		wait for Clk_period;
		Addr <=  "00011000010010";
		Trees_din <= x"1c003a04";
		wait for Clk_period;
		Addr <=  "00011000010011";
		Trees_din <= x"ffd21855";
		wait for Clk_period;
		Addr <=  "00011000010100";
		Trees_din <= x"00151855";
		wait for Clk_period;
		Addr <=  "00011000010101";
		Trees_din <= x"000c100c";
		wait for Clk_period;
		Addr <=  "00011000010110";
		Trees_din <= x"07005404";
		wait for Clk_period;
		Addr <=  "00011000010111";
		Trees_din <= x"00041881";
		wait for Clk_period;
		Addr <=  "00011000011000";
		Trees_din <= x"0c00c904";
		wait for Clk_period;
		Addr <=  "00011000011001";
		Trees_din <= x"ffce1881";
		wait for Clk_period;
		Addr <=  "00011000011010";
		Trees_din <= x"00021881";
		wait for Clk_period;
		Addr <=  "00011000011011";
		Trees_din <= x"07005404";
		wait for Clk_period;
		Addr <=  "00011000011100";
		Trees_din <= x"fff41881";
		wait for Clk_period;
		Addr <=  "00011000011101";
		Trees_din <= x"06fdd504";
		wait for Clk_period;
		Addr <=  "00011000011110";
		Trees_din <= x"002f1881";
		wait for Clk_period;
		Addr <=  "00011000011111";
		Trees_din <= x"00051881";
		wait for Clk_period;
		Addr <=  "00011000100000";
		Trees_din <= x"000e0614";
		wait for Clk_period;
		Addr <=  "00011000100001";
		Trees_din <= x"15faaf04";
		wait for Clk_period;
		Addr <=  "00011000100010";
		Trees_din <= x"ffd518ad";
		wait for Clk_period;
		Addr <=  "00011000100011";
		Trees_din <= x"07005608";
		wait for Clk_period;
		Addr <=  "00011000100100";
		Trees_din <= x"0c00e704";
		wait for Clk_period;
		Addr <=  "00011000100101";
		Trees_din <= x"000518ad";
		wait for Clk_period;
		Addr <=  "00011000100110";
		Trees_din <= x"ffdb18ad";
		wait for Clk_period;
		Addr <=  "00011000100111";
		Trees_din <= x"02012d04";
		wait for Clk_period;
		Addr <=  "00011000101000";
		Trees_din <= x"003318ad";
		wait for Clk_period;
		Addr <=  "00011000101001";
		Trees_din <= x"fff918ad";
		wait for Clk_period;
		Addr <=  "00011000101010";
		Trees_din <= x"001f18ad";
		wait for Clk_period;
		Addr <=  "00011000101011";
		Trees_din <= x"000a0704";
		wait for Clk_period;
		Addr <=  "00011000101100";
		Trees_din <= x"ffe018d1";
		wait for Clk_period;
		Addr <=  "00011000101101";
		Trees_din <= x"11008704";
		wait for Clk_period;
		Addr <=  "00011000101110";
		Trees_din <= x"fff118d1";
		wait for Clk_period;
		Addr <=  "00011000101111";
		Trees_din <= x"15fa8d04";
		wait for Clk_period;
		Addr <=  "00011000110000";
		Trees_din <= x"fff318d1";
		wait for Clk_period;
		Addr <=  "00011000110001";
		Trees_din <= x"0b004204";
		wait for Clk_period;
		Addr <=  "00011000110010";
		Trees_din <= x"000418d1";
		wait for Clk_period;
		Addr <=  "00011000110011";
		Trees_din <= x"003518d1";
		wait for Clk_period;
		Addr <=  "00011000110100";
		Trees_din <= x"1c00380c";
		wait for Clk_period;
		Addr <=  "00011000110101";
		Trees_din <= x"000b6404";
		wait for Clk_period;
		Addr <=  "00011000110110";
		Trees_din <= x"fff118f5";
		wait for Clk_period;
		Addr <=  "00011000110111";
		Trees_din <= x"0f00f504";
		wait for Clk_period;
		Addr <=  "00011000111000";
		Trees_din <= x"000118f5";
		wait for Clk_period;
		Addr <=  "00011000111001";
		Trees_din <= x"003518f5";
		wait for Clk_period;
		Addr <=  "00011000111010";
		Trees_din <= x"04feff04";
		wait for Clk_period;
		Addr <=  "00011000111011";
		Trees_din <= x"ffdb18f5";
		wait for Clk_period;
		Addr <=  "00011000111100";
		Trees_din <= x"000f18f5";
		wait for Clk_period;
		Addr <=  "00011000111101";
		Trees_din <= x"10011b08";
		wait for Clk_period;
		Addr <=  "00011000111110";
		Trees_din <= x"03fcf104";
		wait for Clk_period;
		Addr <=  "00011000111111";
		Trees_din <= x"fff91919";
		wait for Clk_period;
		Addr <=  "00011001000000";
		Trees_din <= x"002a1919";
		wait for Clk_period;
		Addr <=  "00011001000001";
		Trees_din <= x"16007d08";
		wait for Clk_period;
		Addr <=  "00011001000010";
		Trees_din <= x"1c003604";
		wait for Clk_period;
		Addr <=  "00011001000011";
		Trees_din <= x"00081919";
		wait for Clk_period;
		Addr <=  "00011001000100";
		Trees_din <= x"ffd41919";
		wait for Clk_period;
		Addr <=  "00011001000101";
		Trees_din <= x"00101919";
		wait for Clk_period;
		Addr <=  "00011001000110";
		Trees_din <= x"11033710";
		wait for Clk_period;
		Addr <=  "00011001000111";
		Trees_din <= x"11018408";
		wait for Clk_period;
		Addr <=  "00011001001000";
		Trees_din <= x"06fe1f04";
		wait for Clk_period;
		Addr <=  "00011001001001";
		Trees_din <= x"0020193d";
		wait for Clk_period;
		Addr <=  "00011001001010";
		Trees_din <= x"ffe8193d";
		wait for Clk_period;
		Addr <=  "00011001001011";
		Trees_din <= x"0c00c704";
		wait for Clk_period;
		Addr <=  "00011001001100";
		Trees_din <= x"ffd4193d";
		wait for Clk_period;
		Addr <=  "00011001001101";
		Trees_din <= x"0000193d";
		wait for Clk_period;
		Addr <=  "00011001001110";
		Trees_din <= x"001a193d";
		wait for Clk_period;
		Addr <=  "00011001001111";
		Trees_din <= x"10011b08";
		wait for Clk_period;
		Addr <=  "00011001010000";
		Trees_din <= x"03fcf104";
		wait for Clk_period;
		Addr <=  "00011001010001";
		Trees_din <= x"fffb1961";
		wait for Clk_period;
		Addr <=  "00011001010010";
		Trees_din <= x"00261961";
		wait for Clk_period;
		Addr <=  "00011001010011";
		Trees_din <= x"17004708";
		wait for Clk_period;
		Addr <=  "00011001010100";
		Trees_din <= x"18003804";
		wait for Clk_period;
		Addr <=  "00011001010101";
		Trees_din <= x"00091961";
		wait for Clk_period;
		Addr <=  "00011001010110";
		Trees_din <= x"ffcf1961";
		wait for Clk_period;
		Addr <=  "00011001010111";
		Trees_din <= x"00101961";
		wait for Clk_period;
		Addr <=  "00011001011000";
		Trees_din <= x"000b0b08";
		wait for Clk_period;
		Addr <=  "00011001011001";
		Trees_din <= x"12009504";
		wait for Clk_period;
		Addr <=  "00011001011010";
		Trees_din <= x"fffd1985";
		wait for Clk_period;
		Addr <=  "00011001011011";
		Trees_din <= x"ffdb1985";
		wait for Clk_period;
		Addr <=  "00011001011100";
		Trees_din <= x"11008704";
		wait for Clk_period;
		Addr <=  "00011001011101";
		Trees_din <= x"fff11985";
		wait for Clk_period;
		Addr <=  "00011001011110";
		Trees_din <= x"0f00d904";
		wait for Clk_period;
		Addr <=  "00011001011111";
		Trees_din <= x"00031985";
		wait for Clk_period;
		Addr <=  "00011001100000";
		Trees_din <= x"002a1985";
		wait for Clk_period;
		Addr <=  "00011001100001";
		Trees_din <= x"000c100c";
		wait for Clk_period;
		Addr <=  "00011001100010";
		Trees_din <= x"14014c04";
		wait for Clk_period;
		Addr <=  "00011001100011";
		Trees_din <= x"000619b1";
		wait for Clk_period;
		Addr <=  "00011001100100";
		Trees_din <= x"16019d04";
		wait for Clk_period;
		Addr <=  "00011001100101";
		Trees_din <= x"ffd919b1";
		wait for Clk_period;
		Addr <=  "00011001100110";
		Trees_din <= x"fffa19b1";
		wait for Clk_period;
		Addr <=  "00011001100111";
		Trees_din <= x"01fbe308";
		wait for Clk_period;
		Addr <=  "00011001101000";
		Trees_din <= x"19008f04";
		wait for Clk_period;
		Addr <=  "00011001101001";
		Trees_din <= x"ffeb19b1";
		wait for Clk_period;
		Addr <=  "00011001101010";
		Trees_din <= x"001619b1";
		wait for Clk_period;
		Addr <=  "00011001101011";
		Trees_din <= x"002919b1";
		wait for Clk_period;
		Addr <=  "00011001101100";
		Trees_din <= x"11031210";
		wait for Clk_period;
		Addr <=  "00011001101101";
		Trees_din <= x"000e060c";
		wait for Clk_period;
		Addr <=  "00011001101110";
		Trees_din <= x"07005608";
		wait for Clk_period;
		Addr <=  "00011001101111";
		Trees_din <= x"1e005f04";
		wait for Clk_period;
		Addr <=  "00011001110000";
		Trees_din <= x"fff619d5";
		wait for Clk_period;
		Addr <=  "00011001110001";
		Trees_din <= x"ffca19d5";
		wait for Clk_period;
		Addr <=  "00011001110010";
		Trees_din <= x"000c19d5";
		wait for Clk_period;
		Addr <=  "00011001110011";
		Trees_din <= x"001619d5";
		wait for Clk_period;
		Addr <=  "00011001110100";
		Trees_din <= x"001619d5";
		wait for Clk_period;
		Addr <=  "00011001110101";
		Trees_din <= x"15fa8d04";
		wait for Clk_period;
		Addr <=  "00011001110110";
		Trees_din <= x"ffeb19f9";
		wait for Clk_period;
		Addr <=  "00011001110111";
		Trees_din <= x"06ff1b0c";
		wait for Clk_period;
		Addr <=  "00011001111000";
		Trees_din <= x"1504f208";
		wait for Clk_period;
		Addr <=  "00011001111001";
		Trees_din <= x"000bb804";
		wait for Clk_period;
		Addr <=  "00011001111010";
		Trees_din <= x"000019f9";
		wait for Clk_period;
		Addr <=  "00011001111011";
		Trees_din <= x"003019f9";
		wait for Clk_period;
		Addr <=  "00011001111100";
		Trees_din <= x"fff219f9";
		wait for Clk_period;
		Addr <=  "00011001111101";
		Trees_din <= x"ffe819f9";
		wait for Clk_period;
		Addr <=  "00011001111110";
		Trees_din <= x"11033710";
		wait for Clk_period;
		Addr <=  "00011001111111";
		Trees_din <= x"1c002f04";
		wait for Clk_period;
		Addr <=  "00011010000000";
		Trees_din <= x"00131a1d";
		wait for Clk_period;
		Addr <=  "00011010000001";
		Trees_din <= x"0d036408";
		wait for Clk_period;
		Addr <=  "00011010000010";
		Trees_din <= x"1c003a04";
		wait for Clk_period;
		Addr <=  "00011010000011";
		Trees_din <= x"ffcf1a1d";
		wait for Clk_period;
		Addr <=  "00011010000100";
		Trees_din <= x"00041a1d";
		wait for Clk_period;
		Addr <=  "00011010000101";
		Trees_din <= x"00101a1d";
		wait for Clk_period;
		Addr <=  "00011010000110";
		Trees_din <= x"00161a1d";
		wait for Clk_period;
		Addr <=  "00011010000111";
		Trees_din <= x"1c003808";
		wait for Clk_period;
		Addr <=  "00011010001000";
		Trees_din <= x"000b6404";
		wait for Clk_period;
		Addr <=  "00011010001001";
		Trees_din <= x"fff11a39";
		wait for Clk_period;
		Addr <=  "00011010001010";
		Trees_din <= x"00221a39";
		wait for Clk_period;
		Addr <=  "00011010001011";
		Trees_din <= x"04feff04";
		wait for Clk_period;
		Addr <=  "00011010001100";
		Trees_din <= x"ffe11a39";
		wait for Clk_period;
		Addr <=  "00011010001101";
		Trees_din <= x"000a1a39";
		wait for Clk_period;
		Addr <=  "00011010001110";
		Trees_din <= x"11034510";
		wait for Clk_period;
		Addr <=  "00011010001111";
		Trees_din <= x"11018408";
		wait for Clk_period;
		Addr <=  "00011010010000";
		Trees_din <= x"06fe1f04";
		wait for Clk_period;
		Addr <=  "00011010010001";
		Trees_din <= x"001d1a5d";
		wait for Clk_period;
		Addr <=  "00011010010010";
		Trees_din <= x"ffeb1a5d";
		wait for Clk_period;
		Addr <=  "00011010010011";
		Trees_din <= x"02004104";
		wait for Clk_period;
		Addr <=  "00011010010100";
		Trees_din <= x"ffdb1a5d";
		wait for Clk_period;
		Addr <=  "00011010010101";
		Trees_din <= x"00031a5d";
		wait for Clk_period;
		Addr <=  "00011010010110";
		Trees_din <= x"00161a5d";
		wait for Clk_period;
		Addr <=  "00011010010111";
		Trees_din <= x"1c003808";
		wait for Clk_period;
		Addr <=  "00011010011000";
		Trees_din <= x"000b6404";
		wait for Clk_period;
		Addr <=  "00011010011001";
		Trees_din <= x"fff21a79";
		wait for Clk_period;
		Addr <=  "00011010011010";
		Trees_din <= x"00211a79";
		wait for Clk_period;
		Addr <=  "00011010011011";
		Trees_din <= x"06fce904";
		wait for Clk_period;
		Addr <=  "00011010011100";
		Trees_din <= x"ffe01a79";
		wait for Clk_period;
		Addr <=  "00011010011101";
		Trees_din <= x"00061a79";
		wait for Clk_period;
		Addr <=  "00011010011110";
		Trees_din <= x"06ff1b10";
		wait for Clk_period;
		Addr <=  "00011010011111";
		Trees_din <= x"04fecb08";
		wait for Clk_period;
		Addr <=  "00011010100000";
		Trees_din <= x"01fa6c04";
		wait for Clk_period;
		Addr <=  "00011010100001";
		Trees_din <= x"000b1a9d";
		wait for Clk_period;
		Addr <=  "00011010100010";
		Trees_din <= x"ffe41a9d";
		wait for Clk_period;
		Addr <=  "00011010100011";
		Trees_din <= x"0c00c704";
		wait for Clk_period;
		Addr <=  "00011010100100";
		Trees_din <= x"00061a9d";
		wait for Clk_period;
		Addr <=  "00011010100101";
		Trees_din <= x"00281a9d";
		wait for Clk_period;
		Addr <=  "00011010100110";
		Trees_din <= x"ffed1a9d";
		wait for Clk_period;
		Addr <=  "00011010100111";
		Trees_din <= x"10011308";
		wait for Clk_period;
		Addr <=  "00011010101000";
		Trees_din <= x"03fcf104";
		wait for Clk_period;
		Addr <=  "00011010101001";
		Trees_din <= x"fffa1ac1";
		wait for Clk_period;
		Addr <=  "00011010101010";
		Trees_din <= x"00231ac1";
		wait for Clk_period;
		Addr <=  "00011010101011";
		Trees_din <= x"1e006404";
		wait for Clk_period;
		Addr <=  "00011010101100";
		Trees_din <= x"00101ac1";
		wait for Clk_period;
		Addr <=  "00011010101101";
		Trees_din <= x"18003a04";
		wait for Clk_period;
		Addr <=  "00011010101110";
		Trees_din <= x"ffd11ac1";
		wait for Clk_period;
		Addr <=  "00011010101111";
		Trees_din <= x"00051ac1";
		wait for Clk_period;
		Addr <=  "00011010110000";
		Trees_din <= x"0ef96904";
		wait for Clk_period;
		Addr <=  "00011010110001";
		Trees_din <= x"00161ae5";
		wait for Clk_period;
		Addr <=  "00011010110010";
		Trees_din <= x"000e060c";
		wait for Clk_period;
		Addr <=  "00011010110011";
		Trees_din <= x"07005604";
		wait for Clk_period;
		Addr <=  "00011010110100";
		Trees_din <= x"ffda1ae5";
		wait for Clk_period;
		Addr <=  "00011010110101";
		Trees_din <= x"0d01cf04";
		wait for Clk_period;
		Addr <=  "00011010110110";
		Trees_din <= x"00111ae5";
		wait for Clk_period;
		Addr <=  "00011010110111";
		Trees_din <= x"fff71ae5";
		wait for Clk_period;
		Addr <=  "00011010111000";
		Trees_din <= x"001b1ae5";
		wait for Clk_period;
		Addr <=  "00011010111001";
		Trees_din <= x"1c003808";
		wait for Clk_period;
		Addr <=  "00011010111010";
		Trees_din <= x"06fcda04";
		wait for Clk_period;
		Addr <=  "00011010111011";
		Trees_din <= x"00241b01";
		wait for Clk_period;
		Addr <=  "00011010111100";
		Trees_din <= x"fff61b01";
		wait for Clk_period;
		Addr <=  "00011010111101";
		Trees_din <= x"000c1004";
		wait for Clk_period;
		Addr <=  "00011010111110";
		Trees_din <= x"ffe41b01";
		wait for Clk_period;
		Addr <=  "00011010111111";
		Trees_din <= x"00091b01";
		wait for Clk_period;
		Addr <=  "00011011000000";
		Trees_din <= x"15fa8d04";
		wait for Clk_period;
		Addr <=  "00011011000001";
		Trees_din <= x"ffef1b25";
		wait for Clk_period;
		Addr <=  "00011011000010";
		Trees_din <= x"06fed10c";
		wait for Clk_period;
		Addr <=  "00011011000011";
		Trees_din <= x"12008e04";
		wait for Clk_period;
		Addr <=  "00011011000100";
		Trees_din <= x"fff41b25";
		wait for Clk_period;
		Addr <=  "00011011000101";
		Trees_din <= x"16006004";
		wait for Clk_period;
		Addr <=  "00011011000110";
		Trees_din <= x"00361b25";
		wait for Clk_period;
		Addr <=  "00011011000111";
		Trees_din <= x"00001b25";
		wait for Clk_period;
		Addr <=  "00011011001000";
		Trees_din <= x"ffef1b25";
		wait for Clk_period;
		Addr <=  "00011011001001";
		Trees_din <= x"10011308";
		wait for Clk_period;
		Addr <=  "00011011001010";
		Trees_din <= x"1600f104";
		wait for Clk_period;
		Addr <=  "00011011001011";
		Trees_din <= x"001b1b49";
		wait for Clk_period;
		Addr <=  "00011011001100";
		Trees_din <= x"fff81b49";
		wait for Clk_period;
		Addr <=  "00011011001101";
		Trees_din <= x"16007d08";
		wait for Clk_period;
		Addr <=  "00011011001110";
		Trees_din <= x"0f028704";
		wait for Clk_period;
		Addr <=  "00011011001111";
		Trees_din <= x"00011b49";
		wait for Clk_period;
		Addr <=  "00011011010000";
		Trees_din <= x"ffdd1b49";
		wait for Clk_period;
		Addr <=  "00011011010001";
		Trees_din <= x"00101b49";
		wait for Clk_period;
		Addr <=  "00011011010010";
		Trees_din <= x"0a001304";
		wait for Clk_period;
		Addr <=  "00011011010011";
		Trees_din <= x"ffee1b65";
		wait for Clk_period;
		Addr <=  "00011011010100";
		Trees_din <= x"19008f04";
		wait for Clk_period;
		Addr <=  "00011011010101";
		Trees_din <= x"fff01b65";
		wait for Clk_period;
		Addr <=  "00011011010110";
		Trees_din <= x"000b0b04";
		wait for Clk_period;
		Addr <=  "00011011010111";
		Trees_din <= x"fff21b65";
		wait for Clk_period;
		Addr <=  "00011011011000";
		Trees_din <= x"00281b65";
		wait for Clk_period;
		Addr <=  "00011011011001";
		Trees_din <= x"0ef96904";
		wait for Clk_period;
		Addr <=  "00011011011010";
		Trees_din <= x"00131b81";
		wait for Clk_period;
		Addr <=  "00011011011011";
		Trees_din <= x"000e0608";
		wait for Clk_period;
		Addr <=  "00011011011100";
		Trees_din <= x"07005604";
		wait for Clk_period;
		Addr <=  "00011011011101";
		Trees_din <= x"ffdd1b81";
		wait for Clk_period;
		Addr <=  "00011011011110";
		Trees_din <= x"00051b81";
		wait for Clk_period;
		Addr <=  "00011011011111";
		Trees_din <= x"001a1b81";
		wait for Clk_period;
		Addr <=  "00011011100000";
		Trees_din <= x"0effc30c";
		wait for Clk_period;
		Addr <=  "00011011100001";
		Trees_din <= x"0a01f108";
		wait for Clk_period;
		Addr <=  "00011011100010";
		Trees_din <= x"10011304";
		wait for Clk_period;
		Addr <=  "00011011100011";
		Trees_din <= x"00011b9d";
		wait for Clk_period;
		Addr <=  "00011011100100";
		Trees_din <= x"ffd91b9d";
		wait for Clk_period;
		Addr <=  "00011011100101";
		Trees_din <= x"00111b9d";
		wait for Clk_period;
		Addr <=  "00011011100110";
		Trees_din <= x"00111b9d";
		wait for Clk_period;
		Addr <=  "00011011100111";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  2
        -----------
		Addr <=  "00000000000000";
		Trees_din <= x"0610f120";
		wait for Clk_period;
		Addr <=  "00000000000001";
		Trees_din <= x"060d1814";
		wait for Clk_period;
		Addr <=  "00000000000010";
		Trees_din <= x"06088904";
		wait for Clk_period;
		Addr <=  "00000000000011";
		Trees_din <= x"ff4d006d";
		wait for Clk_period;
		Addr <=  "00000000000100";
		Trees_din <= x"00f4590c";
		wait for Clk_period;
		Addr <=  "00000000000101";
		Trees_din <= x"02019008";
		wait for Clk_period;
		Addr <=  "00000000000110";
		Trees_din <= x"02ff7004";
		wait for Clk_period;
		Addr <=  "00000000000111";
		Trees_din <= x"ff78006d";
		wait for Clk_period;
		Addr <=  "00000000001000";
		Trees_din <= x"0187006d";
		wait for Clk_period;
		Addr <=  "00000000001001";
		Trees_din <= x"ff53006d";
		wait for Clk_period;
		Addr <=  "00000000001010";
		Trees_din <= x"02ca006d";
		wait for Clk_period;
		Addr <=  "00000000001011";
		Trees_din <= x"00da7d08";
		wait for Clk_period;
		Addr <=  "00000000001100";
		Trees_din <= x"00ce5b04";
		wait for Clk_period;
		Addr <=  "00000000001101";
		Trees_din <= x"ff59006d";
		wait for Clk_period;
		Addr <=  "00000000001110";
		Trees_din <= x"0027006d";
		wait for Clk_period;
		Addr <=  "00000000001111";
		Trees_din <= x"0383006d";
		wait for Clk_period;
		Addr <=  "00000000010000";
		Trees_din <= x"0211e90c";
		wait for Clk_period;
		Addr <=  "00000000010001";
		Trees_din <= x"011fa004";
		wait for Clk_period;
		Addr <=  "00000000010010";
		Trees_din <= x"041a006d";
		wait for Clk_period;
		Addr <=  "00000000010011";
		Trees_din <= x"03086904";
		wait for Clk_period;
		Addr <=  "00000000010100";
		Trees_din <= x"ff81006d";
		wait for Clk_period;
		Addr <=  "00000000010101";
		Trees_din <= x"00b2006d";
		wait for Clk_period;
		Addr <=  "00000000010110";
		Trees_din <= x"16001708";
		wait for Clk_period;
		Addr <=  "00000000010111";
		Trees_din <= x"05060904";
		wait for Clk_period;
		Addr <=  "00000000011000";
		Trees_din <= x"0027006d";
		wait for Clk_period;
		Addr <=  "00000000011001";
		Trees_din <= x"013c006d";
		wait for Clk_period;
		Addr <=  "00000000011010";
		Trees_din <= x"ff6a006d";
		wait for Clk_period;
		Addr <=  "00000000011011";
		Trees_din <= x"060d1820";
		wait for Clk_period;
		Addr <=  "00000000011100";
		Trees_din <= x"0608890c";
		wait for Clk_period;
		Addr <=  "00000000011101";
		Trees_din <= x"06080304";
		wait for Clk_period;
		Addr <=  "00000000011110";
		Trees_din <= x"ff5400f9";
		wait for Clk_period;
		Addr <=  "00000000011111";
		Trees_din <= x"0ffea004";
		wait for Clk_period;
		Addr <=  "00000000100000";
		Trees_din <= x"004100f9";
		wait for Clk_period;
		Addr <=  "00000000100001";
		Trees_din <= x"ff7100f9";
		wait for Clk_period;
		Addr <=  "00000000100010";
		Trees_din <= x"00ec0008";
		wait for Clk_period;
		Addr <=  "00000000100011";
		Trees_din <= x"1d010c04";
		wait for Clk_period;
		Addr <=  "00000000100100";
		Trees_din <= x"ff5900f9";
		wait for Clk_period;
		Addr <=  "00000000100101";
		Trees_din <= x"003200f9";
		wait for Clk_period;
		Addr <=  "00000000100110";
		Trees_din <= x"13036d08";
		wait for Clk_period;
		Addr <=  "00000000100111";
		Trees_din <= x"02019004";
		wait for Clk_period;
		Addr <=  "00000000101000";
		Trees_din <= x"01cf00f9";
		wait for Clk_period;
		Addr <=  "00000000101001";
		Trees_din <= x"005d00f9";
		wait for Clk_period;
		Addr <=  "00000000101010";
		Trees_din <= x"ff9d00f9";
		wait for Clk_period;
		Addr <=  "00000000101011";
		Trees_din <= x"02145120";
		wait for Clk_period;
		Addr <=  "00000000101100";
		Trees_din <= x"011cba14";
		wait for Clk_period;
		Addr <=  "00000000101101";
		Trees_din <= x"0312d510";
		wait for Clk_period;
		Addr <=  "00000000101110";
		Trees_din <= x"05098d08";
		wait for Clk_period;
		Addr <=  "00000000101111";
		Trees_din <= x"04171604";
		wait for Clk_period;
		Addr <=  "00000000110000";
		Trees_din <= x"01b000f9";
		wait for Clk_period;
		Addr <=  "00000000110001";
		Trees_din <= x"00ad00f9";
		wait for Clk_period;
		Addr <=  "00000000110010";
		Trees_din <= x"0a006104";
		wait for Clk_period;
		Addr <=  "00000000110011";
		Trees_din <= x"00b200f9";
		wait for Clk_period;
		Addr <=  "00000000110100";
		Trees_din <= x"003000f9";
		wait for Clk_period;
		Addr <=  "00000000110101";
		Trees_din <= x"ff9700f9";
		wait for Clk_period;
		Addr <=  "00000000110110";
		Trees_din <= x"0615fc04";
		wait for Clk_period;
		Addr <=  "00000000110111";
		Trees_din <= x"ff6200f9";
		wait for Clk_period;
		Addr <=  "00000000111000";
		Trees_din <= x"15027e04";
		wait for Clk_period;
		Addr <=  "00000000111001";
		Trees_din <= x"019b00f9";
		wait for Clk_period;
		Addr <=  "00000000111010";
		Trees_din <= x"002500f9";
		wait for Clk_period;
		Addr <=  "00000000111011";
		Trees_din <= x"1f040004";
		wait for Clk_period;
		Addr <=  "00000000111100";
		Trees_din <= x"002900f9";
		wait for Clk_period;
		Addr <=  "00000000111101";
		Trees_din <= x"ff6400f9";
		wait for Clk_period;
		Addr <=  "00000000111110";
		Trees_din <= x"060d1820";
		wait for Clk_period;
		Addr <=  "00000000111111";
		Trees_din <= x"0608890c";
		wait for Clk_period;
		Addr <=  "00000001000000";
		Trees_din <= x"0e059f04";
		wait for Clk_period;
		Addr <=  "00000001000001";
		Trees_din <= x"ff59017d";
		wait for Clk_period;
		Addr <=  "00000001000010";
		Trees_din <= x"0d00f204";
		wait for Clk_period;
		Addr <=  "00000001000011";
		Trees_din <= x"003e017d";
		wait for Clk_period;
		Addr <=  "00000001000100";
		Trees_din <= x"ff7b017d";
		wait for Clk_period;
		Addr <=  "00000001000101";
		Trees_din <= x"00ec0008";
		wait for Clk_period;
		Addr <=  "00000001000110";
		Trees_din <= x"1d010c04";
		wait for Clk_period;
		Addr <=  "00000001000111";
		Trees_din <= x"ff5f017d";
		wait for Clk_period;
		Addr <=  "00000001001000";
		Trees_din <= x"002f017d";
		wait for Clk_period;
		Addr <=  "00000001001001";
		Trees_din <= x"01fb0804";
		wait for Clk_period;
		Addr <=  "00000001001010";
		Trees_din <= x"fffa017d";
		wait for Clk_period;
		Addr <=  "00000001001011";
		Trees_din <= x"0b026504";
		wait for Clk_period;
		Addr <=  "00000001001100";
		Trees_din <= x"0132017d";
		wait for Clk_period;
		Addr <=  "00000001001101";
		Trees_din <= x"001d017d";
		wait for Clk_period;
		Addr <=  "00000001001110";
		Trees_din <= x"0214511c";
		wait for Clk_period;
		Addr <=  "00000001001111";
		Trees_din <= x"011fa014";
		wait for Clk_period;
		Addr <=  "00000001010000";
		Trees_din <= x"050bc110";
		wait for Clk_period;
		Addr <=  "00000001010001";
		Trees_din <= x"060e1c08";
		wait for Clk_period;
		Addr <=  "00000001010010";
		Trees_din <= x"04015904";
		wait for Clk_period;
		Addr <=  "00000001010011";
		Trees_din <= x"0115017d";
		wait for Clk_period;
		Addr <=  "00000001010100";
		Trees_din <= x"ffbf017d";
		wait for Clk_period;
		Addr <=  "00000001010101";
		Trees_din <= x"01f42104";
		wait for Clk_period;
		Addr <=  "00000001010110";
		Trees_din <= x"005f017d";
		wait for Clk_period;
		Addr <=  "00000001010111";
		Trees_din <= x"0134017d";
		wait for Clk_period;
		Addr <=  "00000001011000";
		Trees_din <= x"ff9b017d";
		wait for Clk_period;
		Addr <=  "00000001011001";
		Trees_din <= x"061cb504";
		wait for Clk_period;
		Addr <=  "00000001011010";
		Trees_din <= x"ff6d017d";
		wait for Clk_period;
		Addr <=  "00000001011011";
		Trees_din <= x"012d017d";
		wait for Clk_period;
		Addr <=  "00000001011100";
		Trees_din <= x"1f040004";
		wait for Clk_period;
		Addr <=  "00000001011101";
		Trees_din <= x"0039017d";
		wait for Clk_period;
		Addr <=  "00000001011110";
		Trees_din <= x"ff6a017d";
		wait for Clk_period;
		Addr <=  "00000001011111";
		Trees_din <= x"060d181c";
		wait for Clk_period;
		Addr <=  "00000001100000";
		Trees_din <= x"06080304";
		wait for Clk_period;
		Addr <=  "00000001100001";
		Trees_din <= x"ff5c01f9";
		wait for Clk_period;
		Addr <=  "00000001100010";
		Trees_din <= x"00ec0008";
		wait for Clk_period;
		Addr <=  "00000001100011";
		Trees_din <= x"1d010c04";
		wait for Clk_period;
		Addr <=  "00000001100100";
		Trees_din <= x"ff6201f9";
		wait for Clk_period;
		Addr <=  "00000001100101";
		Trees_din <= x"002c01f9";
		wait for Clk_period;
		Addr <=  "00000001100110";
		Trees_din <= x"0207240c";
		wait for Clk_period;
		Addr <=  "00000001100111";
		Trees_din <= x"10003304";
		wait for Clk_period;
		Addr <=  "00000001101000";
		Trees_din <= x"002201f9";
		wait for Clk_period;
		Addr <=  "00000001101001";
		Trees_din <= x"05f69a04";
		wait for Clk_period;
		Addr <=  "00000001101010";
		Trees_din <= x"002401f9";
		wait for Clk_period;
		Addr <=  "00000001101011";
		Trees_din <= x"012101f9";
		wait for Clk_period;
		Addr <=  "00000001101100";
		Trees_din <= x"ffa701f9";
		wait for Clk_period;
		Addr <=  "00000001101101";
		Trees_din <= x"0214511c";
		wait for Clk_period;
		Addr <=  "00000001101110";
		Trees_din <= x"011fa014";
		wait for Clk_period;
		Addr <=  "00000001101111";
		Trees_din <= x"050bc110";
		wait for Clk_period;
		Addr <=  "00000001110000";
		Trees_din <= x"060f9508";
		wait for Clk_period;
		Addr <=  "00000001110001";
		Trees_din <= x"01081b04";
		wait for Clk_period;
		Addr <=  "00000001110010";
		Trees_din <= x"00e501f9";
		wait for Clk_period;
		Addr <=  "00000001110011";
		Trees_din <= x"ff8301f9";
		wait for Clk_period;
		Addr <=  "00000001110100";
		Trees_din <= x"01f42104";
		wait for Clk_period;
		Addr <=  "00000001110101";
		Trees_din <= x"004f01f9";
		wait for Clk_period;
		Addr <=  "00000001110110";
		Trees_din <= x"00fc01f9";
		wait for Clk_period;
		Addr <=  "00000001110111";
		Trees_din <= x"ffa401f9";
		wait for Clk_period;
		Addr <=  "00000001111000";
		Trees_din <= x"061cb504";
		wait for Clk_period;
		Addr <=  "00000001111001";
		Trees_din <= x"ff7401f9";
		wait for Clk_period;
		Addr <=  "00000001111010";
		Trees_din <= x"00f001f9";
		wait for Clk_period;
		Addr <=  "00000001111011";
		Trees_din <= x"0a02ce04";
		wait for Clk_period;
		Addr <=  "00000001111100";
		Trees_din <= x"ff6f01f9";
		wait for Clk_period;
		Addr <=  "00000001111101";
		Trees_din <= x"003801f9";
		wait for Clk_period;
		Addr <=  "00000001111110";
		Trees_din <= x"060af018";
		wait for Clk_period;
		Addr <=  "00000001111111";
		Trees_din <= x"06080304";
		wait for Clk_period;
		Addr <=  "00000010000000";
		Trees_din <= x"ff5f0275";
		wait for Clk_period;
		Addr <=  "00000010000001";
		Trees_din <= x"00f4590c";
		wait for Clk_period;
		Addr <=  "00000010000010";
		Trees_din <= x"10034504";
		wait for Clk_period;
		Addr <=  "00000010000011";
		Trees_din <= x"ff6a0275";
		wait for Clk_period;
		Addr <=  "00000010000100";
		Trees_din <= x"0200d404";
		wait for Clk_period;
		Addr <=  "00000010000101";
		Trees_din <= x"007a0275";
		wait for Clk_period;
		Addr <=  "00000010000110";
		Trees_din <= x"ffa00275";
		wait for Clk_period;
		Addr <=  "00000010000111";
		Trees_din <= x"10001904";
		wait for Clk_period;
		Addr <=  "00000010001000";
		Trees_din <= x"00100275";
		wait for Clk_period;
		Addr <=  "00000010001001";
		Trees_din <= x"00dc0275";
		wait for Clk_period;
		Addr <=  "00000010001010";
		Trees_din <= x"02145120";
		wait for Clk_period;
		Addr <=  "00000010001011";
		Trees_din <= x"011cba14";
		wait for Clk_period;
		Addr <=  "00000010001100";
		Trees_din <= x"0312d510";
		wait for Clk_period;
		Addr <=  "00000010001101";
		Trees_din <= x"060e1c08";
		wait for Clk_period;
		Addr <=  "00000010001110";
		Trees_din <= x"00da7d04";
		wait for Clk_period;
		Addr <=  "00000010001111";
		Trees_din <= x"ff830275";
		wait for Clk_period;
		Addr <=  "00000010010000";
		Trees_din <= x"00c50275";
		wait for Clk_period;
		Addr <=  "00000010010001";
		Trees_din <= x"04171604";
		wait for Clk_period;
		Addr <=  "00000010010010";
		Trees_din <= x"00dc0275";
		wait for Clk_period;
		Addr <=  "00000010010011";
		Trees_din <= x"00630275";
		wait for Clk_period;
		Addr <=  "00000010010100";
		Trees_din <= x"ff8f0275";
		wait for Clk_period;
		Addr <=  "00000010010101";
		Trees_din <= x"0615fc04";
		wait for Clk_period;
		Addr <=  "00000010010110";
		Trees_din <= x"ff720275";
		wait for Clk_period;
		Addr <=  "00000010010111";
		Trees_din <= x"15027e04";
		wait for Clk_period;
		Addr <=  "00000010011000";
		Trees_din <= x"00d30275";
		wait for Clk_period;
		Addr <=  "00000010011001";
		Trees_din <= x"00120275";
		wait for Clk_period;
		Addr <=  "00000010011010";
		Trees_din <= x"0a03ba04";
		wait for Clk_period;
		Addr <=  "00000010011011";
		Trees_din <= x"ff6e0275";
		wait for Clk_period;
		Addr <=  "00000010011100";
		Trees_din <= x"00390275";
		wait for Clk_period;
		Addr <=  "00000010011101";
		Trees_din <= x"060af014";
		wait for Clk_period;
		Addr <=  "00000010011110";
		Trees_din <= x"06080304";
		wait for Clk_period;
		Addr <=  "00000010011111";
		Trees_din <= x"ff6102e9";
		wait for Clk_period;
		Addr <=  "00000010100000";
		Trees_din <= x"00ecda04";
		wait for Clk_period;
		Addr <=  "00000010100001";
		Trees_din <= x"ff7002e9";
		wait for Clk_period;
		Addr <=  "00000010100010";
		Trees_din <= x"05fc1404";
		wait for Clk_period;
		Addr <=  "00000010100011";
		Trees_din <= x"ffd602e9";
		wait for Clk_period;
		Addr <=  "00000010100100";
		Trees_din <= x"09043d04";
		wait for Clk_period;
		Addr <=  "00000010100101";
		Trees_din <= x"00c102e9";
		wait for Clk_period;
		Addr <=  "00000010100110";
		Trees_din <= x"003c02e9";
		wait for Clk_period;
		Addr <=  "00000010100111";
		Trees_din <= x"02145120";
		wait for Clk_period;
		Addr <=  "00000010101000";
		Trees_din <= x"011cba14";
		wait for Clk_period;
		Addr <=  "00000010101001";
		Trees_din <= x"0312d510";
		wait for Clk_period;
		Addr <=  "00000010101010";
		Trees_din <= x"060e1c08";
		wait for Clk_period;
		Addr <=  "00000010101011";
		Trees_din <= x"00da7d04";
		wait for Clk_period;
		Addr <=  "00000010101100";
		Trees_din <= x"ff8b02e9";
		wait for Clk_period;
		Addr <=  "00000010101101";
		Trees_din <= x"00a702e9";
		wait for Clk_period;
		Addr <=  "00000010101110";
		Trees_din <= x"04171604";
		wait for Clk_period;
		Addr <=  "00000010101111";
		Trees_din <= x"00c702e9";
		wait for Clk_period;
		Addr <=  "00000010110000";
		Trees_din <= x"005302e9";
		wait for Clk_period;
		Addr <=  "00000010110001";
		Trees_din <= x"ff9a02e9";
		wait for Clk_period;
		Addr <=  "00000010110010";
		Trees_din <= x"0615fc04";
		wait for Clk_period;
		Addr <=  "00000010110011";
		Trees_din <= x"ff7902e9";
		wait for Clk_period;
		Addr <=  "00000010110100";
		Trees_din <= x"061cb504";
		wait for Clk_period;
		Addr <=  "00000010110101";
		Trees_din <= x"003302e9";
		wait for Clk_period;
		Addr <=  "00000010110110";
		Trees_din <= x"00b402e9";
		wait for Clk_period;
		Addr <=  "00000010110111";
		Trees_din <= x"0a03ba04";
		wait for Clk_period;
		Addr <=  "00000010111000";
		Trees_din <= x"ff7402e9";
		wait for Clk_period;
		Addr <=  "00000010111001";
		Trees_din <= x"003502e9";
		wait for Clk_period;
		Addr <=  "00000010111010";
		Trees_din <= x"060af018";
		wait for Clk_period;
		Addr <=  "00000010111011";
		Trees_din <= x"0608030c";
		wait for Clk_period;
		Addr <=  "00000010111100";
		Trees_din <= x"11000008";
		wait for Clk_period;
		Addr <=  "00000010111101";
		Trees_din <= x"1200a204";
		wait for Clk_period;
		Addr <=  "00000010111110";
		Trees_din <= x"ff7a035d";
		wait for Clk_period;
		Addr <=  "00000010111111";
		Trees_din <= x"003f035d";
		wait for Clk_period;
		Addr <=  "00000011000000";
		Trees_din <= x"ff62035d";
		wait for Clk_period;
		Addr <=  "00000011000001";
		Trees_din <= x"00ecda04";
		wait for Clk_period;
		Addr <=  "00000011000010";
		Trees_din <= x"ff75035d";
		wait for Clk_period;
		Addr <=  "00000011000011";
		Trees_din <= x"05fc1404";
		wait for Clk_period;
		Addr <=  "00000011000100";
		Trees_din <= x"ffdb035d";
		wait for Clk_period;
		Addr <=  "00000011000101";
		Trees_din <= x"0097035d";
		wait for Clk_period;
		Addr <=  "00000011000110";
		Trees_din <= x"0214511c";
		wait for Clk_period;
		Addr <=  "00000011000111";
		Trees_din <= x"011fa014";
		wait for Clk_period;
		Addr <=  "00000011001000";
		Trees_din <= x"050bc110";
		wait for Clk_period;
		Addr <=  "00000011001001";
		Trees_din <= x"060f9508";
		wait for Clk_period;
		Addr <=  "00000011001010";
		Trees_din <= x"00da7d04";
		wait for Clk_period;
		Addr <=  "00000011001011";
		Trees_din <= x"ff8b035d";
		wait for Clk_period;
		Addr <=  "00000011001100";
		Trees_din <= x"0095035d";
		wait for Clk_period;
		Addr <=  "00000011001101";
		Trees_din <= x"01f42104";
		wait for Clk_period;
		Addr <=  "00000011001110";
		Trees_din <= x"002b035d";
		wait for Clk_period;
		Addr <=  "00000011001111";
		Trees_din <= x"00b8035d";
		wait for Clk_period;
		Addr <=  "00000011010000";
		Trees_din <= x"ffa7035d";
		wait for Clk_period;
		Addr <=  "00000011010001";
		Trees_din <= x"061cb504";
		wait for Clk_period;
		Addr <=  "00000011010010";
		Trees_din <= x"ff85035d";
		wait for Clk_period;
		Addr <=  "00000011010011";
		Trees_din <= x"0094035d";
		wait for Clk_period;
		Addr <=  "00000011010100";
		Trees_din <= x"0e015504";
		wait for Clk_period;
		Addr <=  "00000011010101";
		Trees_din <= x"ff7b035d";
		wait for Clk_period;
		Addr <=  "00000011010110";
		Trees_din <= x"0029035d";
		wait for Clk_period;
		Addr <=  "00000011010111";
		Trees_din <= x"060af01c";
		wait for Clk_period;
		Addr <=  "00000011011000";
		Trees_din <= x"0608030c";
		wait for Clk_period;
		Addr <=  "00000011011001";
		Trees_din <= x"11000008";
		wait for Clk_period;
		Addr <=  "00000011011010";
		Trees_din <= x"18003204";
		wait for Clk_period;
		Addr <=  "00000011011011";
		Trees_din <= x"004303e9";
		wait for Clk_period;
		Addr <=  "00000011011100";
		Trees_din <= x"ff8103e9";
		wait for Clk_period;
		Addr <=  "00000011011101";
		Trees_din <= x"ff6303e9";
		wait for Clk_period;
		Addr <=  "00000011011110";
		Trees_din <= x"00ecda04";
		wait for Clk_period;
		Addr <=  "00000011011111";
		Trees_din <= x"ff7b03e9";
		wait for Clk_period;
		Addr <=  "00000011100000";
		Trees_din <= x"05fc1404";
		wait for Clk_period;
		Addr <=  "00000011100001";
		Trees_din <= x"ffe103e9";
		wait for Clk_period;
		Addr <=  "00000011100010";
		Trees_din <= x"09043d04";
		wait for Clk_period;
		Addr <=  "00000011100011";
		Trees_din <= x"009503e9";
		wait for Clk_period;
		Addr <=  "00000011100100";
		Trees_din <= x"002603e9";
		wait for Clk_period;
		Addr <=  "00000011100101";
		Trees_din <= x"02145124";
		wait for Clk_period;
		Addr <=  "00000011100110";
		Trees_din <= x"011cba18";
		wait for Clk_period;
		Addr <=  "00000011100111";
		Trees_din <= x"060e1c0c";
		wait for Clk_period;
		Addr <=  "00000011101000";
		Trees_din <= x"04033104";
		wait for Clk_period;
		Addr <=  "00000011101001";
		Trees_din <= x"009703e9";
		wait for Clk_period;
		Addr <=  "00000011101010";
		Trees_din <= x"0f004a04";
		wait for Clk_period;
		Addr <=  "00000011101011";
		Trees_din <= x"003703e9";
		wait for Clk_period;
		Addr <=  "00000011101100";
		Trees_din <= x"ff7b03e9";
		wait for Clk_period;
		Addr <=  "00000011101101";
		Trees_din <= x"04171608";
		wait for Clk_period;
		Addr <=  "00000011101110";
		Trees_din <= x"07005c04";
		wait for Clk_period;
		Addr <=  "00000011101111";
		Trees_din <= x"00af03e9";
		wait for Clk_period;
		Addr <=  "00000011110000";
		Trees_din <= x"005a03e9";
		wait for Clk_period;
		Addr <=  "00000011110001";
		Trees_din <= x"003103e9";
		wait for Clk_period;
		Addr <=  "00000011110010";
		Trees_din <= x"0615fc04";
		wait for Clk_period;
		Addr <=  "00000011110011";
		Trees_din <= x"ff8703e9";
		wait for Clk_period;
		Addr <=  "00000011110100";
		Trees_din <= x"061cb504";
		wait for Clk_period;
		Addr <=  "00000011110101";
		Trees_din <= x"002a03e9";
		wait for Clk_period;
		Addr <=  "00000011110110";
		Trees_din <= x"008d03e9";
		wait for Clk_period;
		Addr <=  "00000011110111";
		Trees_din <= x"1f040004";
		wait for Clk_period;
		Addr <=  "00000011111000";
		Trees_din <= x"002903e9";
		wait for Clk_period;
		Addr <=  "00000011111001";
		Trees_din <= x"ff8203e9";
		wait for Clk_period;
		Addr <=  "00000011111010";
		Trees_din <= x"06093514";
		wait for Clk_period;
		Addr <=  "00000011111011";
		Trees_din <= x"0608030c";
		wait for Clk_period;
		Addr <=  "00000011111100";
		Trees_din <= x"11000008";
		wait for Clk_period;
		Addr <=  "00000011111101";
		Trees_din <= x"1200a204";
		wait for Clk_period;
		Addr <=  "00000011111110";
		Trees_din <= x"ff87045d";
		wait for Clk_period;
		Addr <=  "00000011111111";
		Trees_din <= x"0044045d";
		wait for Clk_period;
		Addr <=  "00000100000000";
		Trees_din <= x"ff64045d";
		wait for Clk_period;
		Addr <=  "00000100000001";
		Trees_din <= x"00f45904";
		wait for Clk_period;
		Addr <=  "00000100000010";
		Trees_din <= x"ff8b045d";
		wait for Clk_period;
		Addr <=  "00000100000011";
		Trees_din <= x"0060045d";
		wait for Clk_period;
		Addr <=  "00000100000100";
		Trees_din <= x"02145120";
		wait for Clk_period;
		Addr <=  "00000100000101";
		Trees_din <= x"060f9510";
		wait for Clk_period;
		Addr <=  "00000100000110";
		Trees_din <= x"00da7d04";
		wait for Clk_period;
		Addr <=  "00000100000111";
		Trees_din <= x"ff81045d";
		wait for Clk_period;
		Addr <=  "00000100001000";
		Trees_din <= x"02fc1404";
		wait for Clk_period;
		Addr <=  "00000100001001";
		Trees_din <= x"ffdf045d";
		wait for Clk_period;
		Addr <=  "00000100001010";
		Trees_din <= x"02022704";
		wait for Clk_period;
		Addr <=  "00000100001011";
		Trees_din <= x"009d045d";
		wait for Clk_period;
		Addr <=  "00000100001100";
		Trees_din <= x"001d045d";
		wait for Clk_period;
		Addr <=  "00000100001101";
		Trees_din <= x"0123d70c";
		wait for Clk_period;
		Addr <=  "00000100001110";
		Trees_din <= x"04171608";
		wait for Clk_period;
		Addr <=  "00000100001111";
		Trees_din <= x"01f88a04";
		wait for Clk_period;
		Addr <=  "00000100010000";
		Trees_din <= x"0042045d";
		wait for Clk_period;
		Addr <=  "00000100010001";
		Trees_din <= x"00a8045d";
		wait for Clk_period;
		Addr <=  "00000100010010";
		Trees_din <= x"0026045d";
		wait for Clk_period;
		Addr <=  "00000100010011";
		Trees_din <= x"ffe4045d";
		wait for Clk_period;
		Addr <=  "00000100010100";
		Trees_din <= x"0ffea804";
		wait for Clk_period;
		Addr <=  "00000100010101";
		Trees_din <= x"0024045d";
		wait for Clk_period;
		Addr <=  "00000100010110";
		Trees_din <= x"ff80045d";
		wait for Clk_period;
		Addr <=  "00000100010111";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00000100011000";
		Trees_din <= x"060af018";
		wait for Clk_period;
		Addr <=  "00000100011001";
		Trees_din <= x"0608030c";
		wait for Clk_period;
		Addr <=  "00000100011010";
		Trees_din <= x"11000008";
		wait for Clk_period;
		Addr <=  "00000100011011";
		Trees_din <= x"06002c04";
		wait for Clk_period;
		Addr <=  "00000100011100";
		Trees_din <= x"ff8e04d5";
		wait for Clk_period;
		Addr <=  "00000100011101";
		Trees_din <= x"004304d5";
		wait for Clk_period;
		Addr <=  "00000100011110";
		Trees_din <= x"ff6504d5";
		wait for Clk_period;
		Addr <=  "00000100011111";
		Trees_din <= x"00ecda04";
		wait for Clk_period;
		Addr <=  "00000100100000";
		Trees_din <= x"ff8804d5";
		wait for Clk_period;
		Addr <=  "00000100100001";
		Trees_din <= x"05fc1404";
		wait for Clk_period;
		Addr <=  "00000100100010";
		Trees_din <= x"ffe404d5";
		wait for Clk_period;
		Addr <=  "00000100100011";
		Trees_din <= x"006b04d5";
		wait for Clk_period;
		Addr <=  "00000100100100";
		Trees_din <= x"0214511c";
		wait for Clk_period;
		Addr <=  "00000100100101";
		Trees_din <= x"06138014";
		wait for Clk_period;
		Addr <=  "00000100100110";
		Trees_din <= x"00d25d08";
		wait for Clk_period;
		Addr <=  "00000100100111";
		Trees_din <= x"0effeb04";
		wait for Clk_period;
		Addr <=  "00000100101000";
		Trees_din <= x"ff7904d5";
		wait for Clk_period;
		Addr <=  "00000100101001";
		Trees_din <= x"ffeb04d5";
		wait for Clk_period;
		Addr <=  "00000100101010";
		Trees_din <= x"02fa4c04";
		wait for Clk_period;
		Addr <=  "00000100101011";
		Trees_din <= x"ffde04d5";
		wait for Clk_period;
		Addr <=  "00000100101100";
		Trees_din <= x"02063904";
		wait for Clk_period;
		Addr <=  "00000100101101";
		Trees_din <= x"009804d5";
		wait for Clk_period;
		Addr <=  "00000100101110";
		Trees_din <= x"003104d5";
		wait for Clk_period;
		Addr <=  "00000100101111";
		Trees_din <= x"0123d704";
		wait for Clk_period;
		Addr <=  "00000100110000";
		Trees_din <= x"00a504d5";
		wait for Clk_period;
		Addr <=  "00000100110001";
		Trees_din <= x"000204d5";
		wait for Clk_period;
		Addr <=  "00000100110010";
		Trees_din <= x"1100a704";
		wait for Clk_period;
		Addr <=  "00000100110011";
		Trees_din <= x"002204d5";
		wait for Clk_period;
		Addr <=  "00000100110100";
		Trees_din <= x"ff9004d5";
		wait for Clk_period;
		Addr <=  "00000100110101";
		Trees_din <= x"0609350c";
		wait for Clk_period;
		Addr <=  "00000100110110";
		Trees_din <= x"06047104";
		wait for Clk_period;
		Addr <=  "00000100110111";
		Trees_din <= x"ff660529";
		wait for Clk_period;
		Addr <=  "00000100111000";
		Trees_din <= x"00fcab04";
		wait for Clk_period;
		Addr <=  "00000100111001";
		Trees_din <= x"ff830529";
		wait for Clk_period;
		Addr <=  "00000100111010";
		Trees_din <= x"007e0529";
		wait for Clk_period;
		Addr <=  "00000100111011";
		Trees_din <= x"06138018";
		wait for Clk_period;
		Addr <=  "00000100111100";
		Trees_din <= x"00d90008";
		wait for Clk_period;
		Addr <=  "00000100111101";
		Trees_din <= x"05fcf104";
		wait for Clk_period;
		Addr <=  "00000100111110";
		Trees_din <= x"00020529";
		wait for Clk_period;
		Addr <=  "00000100111111";
		Trees_din <= x"ff780529";
		wait for Clk_period;
		Addr <=  "00000101000000";
		Trees_din <= x"02fa4c04";
		wait for Clk_period;
		Addr <=  "00000101000001";
		Trees_din <= x"ffe10529";
		wait for Clk_period;
		Addr <=  "00000101000010";
		Trees_din <= x"02063908";
		wait for Clk_period;
		Addr <=  "00000101000011";
		Trees_din <= x"0c024004";
		wait for Clk_period;
		Addr <=  "00000101000100";
		Trees_din <= x"00940529";
		wait for Clk_period;
		Addr <=  "00000101000101";
		Trees_din <= x"00200529";
		wait for Clk_period;
		Addr <=  "00000101000110";
		Trees_din <= x"001d0529";
		wait for Clk_period;
		Addr <=  "00000101000111";
		Trees_din <= x"0123d704";
		wait for Clk_period;
		Addr <=  "00000101001000";
		Trees_din <= x"009e0529";
		wait for Clk_period;
		Addr <=  "00000101001001";
		Trees_din <= x"ffef0529";
		wait for Clk_period;
		Addr <=  "00000101001010";
		Trees_din <= x"0609350c";
		wait for Clk_period;
		Addr <=  "00000101001011";
		Trees_din <= x"06047104";
		wait for Clk_period;
		Addr <=  "00000101001100";
		Trees_din <= x"ff67058d";
		wait for Clk_period;
		Addr <=  "00000101001101";
		Trees_din <= x"04ff8e04";
		wait for Clk_period;
		Addr <=  "00000101001110";
		Trees_din <= x"0068058d";
		wait for Clk_period;
		Addr <=  "00000101001111";
		Trees_din <= x"ff8a058d";
		wait for Clk_period;
		Addr <=  "00000101010000";
		Trees_din <= x"0610f114";
		wait for Clk_period;
		Addr <=  "00000101010001";
		Trees_din <= x"00ddf608";
		wait for Clk_period;
		Addr <=  "00000101010010";
		Trees_din <= x"0effeb04";
		wait for Clk_period;
		Addr <=  "00000101010011";
		Trees_din <= x"ff86058d";
		wait for Clk_period;
		Addr <=  "00000101010100";
		Trees_din <= x"fff2058d";
		wait for Clk_period;
		Addr <=  "00000101010101";
		Trees_din <= x"0b025f08";
		wait for Clk_period;
		Addr <=  "00000101010110";
		Trees_din <= x"01fc7d04";
		wait for Clk_period;
		Addr <=  "00000101010111";
		Trees_din <= x"0024058d";
		wait for Clk_period;
		Addr <=  "00000101011000";
		Trees_din <= x"0084058d";
		wait for Clk_period;
		Addr <=  "00000101011001";
		Trees_din <= x"ffe0058d";
		wait for Clk_period;
		Addr <=  "00000101011010";
		Trees_din <= x"0123d710";
		wait for Clk_period;
		Addr <=  "00000101011011";
		Trees_din <= x"0417160c";
		wait for Clk_period;
		Addr <=  "00000101011100";
		Trees_din <= x"07005c04";
		wait for Clk_period;
		Addr <=  "00000101011101";
		Trees_din <= x"009a058d";
		wait for Clk_period;
		Addr <=  "00000101011110";
		Trees_din <= x"0615fc04";
		wait for Clk_period;
		Addr <=  "00000101011111";
		Trees_din <= x"fff6058d";
		wait for Clk_period;
		Addr <=  "00000101100000";
		Trees_din <= x"0059058d";
		wait for Clk_period;
		Addr <=  "00000101100001";
		Trees_din <= x"000b058d";
		wait for Clk_period;
		Addr <=  "00000101100010";
		Trees_din <= x"ffe6058d";
		wait for Clk_period;
		Addr <=  "00000101100011";
		Trees_din <= x"0609350c";
		wait for Clk_period;
		Addr <=  "00000101100100";
		Trees_din <= x"06047104";
		wait for Clk_period;
		Addr <=  "00000101100101";
		Trees_din <= x"ff6705e1";
		wait for Clk_period;
		Addr <=  "00000101100110";
		Trees_din <= x"01fe7d04";
		wait for Clk_period;
		Addr <=  "00000101100111";
		Trees_din <= x"004f05e1";
		wait for Clk_period;
		Addr <=  "00000101101000";
		Trees_din <= x"ff8505e1";
		wait for Clk_period;
		Addr <=  "00000101101001";
		Trees_din <= x"06138018";
		wait for Clk_period;
		Addr <=  "00000101101010";
		Trees_din <= x"00d71808";
		wait for Clk_period;
		Addr <=  "00000101101011";
		Trees_din <= x"03018d04";
		wait for Clk_period;
		Addr <=  "00000101101100";
		Trees_din <= x"ffe505e1";
		wait for Clk_period;
		Addr <=  "00000101101101";
		Trees_din <= x"ff8205e1";
		wait for Clk_period;
		Addr <=  "00000101101110";
		Trees_din <= x"02fa4c04";
		wait for Clk_period;
		Addr <=  "00000101101111";
		Trees_din <= x"ffce05e1";
		wait for Clk_period;
		Addr <=  "00000101110000";
		Trees_din <= x"02063908";
		wait for Clk_period;
		Addr <=  "00000101110001";
		Trees_din <= x"0f02a504";
		wait for Clk_period;
		Addr <=  "00000101110010";
		Trees_din <= x"008b05e1";
		wait for Clk_period;
		Addr <=  "00000101110011";
		Trees_din <= x"003005e1";
		wait for Clk_period;
		Addr <=  "00000101110100";
		Trees_din <= x"000e05e1";
		wait for Clk_period;
		Addr <=  "00000101110101";
		Trees_din <= x"0123d704";
		wait for Clk_period;
		Addr <=  "00000101110110";
		Trees_din <= x"009605e1";
		wait for Clk_period;
		Addr <=  "00000101110111";
		Trees_din <= x"fff905e1";
		wait for Clk_period;
		Addr <=  "00000101111000";
		Trees_din <= x"060af010";
		wait for Clk_period;
		Addr <=  "00000101111001";
		Trees_din <= x"06047104";
		wait for Clk_period;
		Addr <=  "00000101111010";
		Trees_din <= x"ff68062d";
		wait for Clk_period;
		Addr <=  "00000101111011";
		Trees_din <= x"00fcab08";
		wait for Clk_period;
		Addr <=  "00000101111100";
		Trees_din <= x"14004604";
		wait for Clk_period;
		Addr <=  "00000101111101";
		Trees_din <= x"ffee062d";
		wait for Clk_period;
		Addr <=  "00000101111110";
		Trees_din <= x"ff8c062d";
		wait for Clk_period;
		Addr <=  "00000101111111";
		Trees_din <= x"006a062d";
		wait for Clk_period;
		Addr <=  "00000110000000";
		Trees_din <= x"06138010";
		wait for Clk_period;
		Addr <=  "00000110000001";
		Trees_din <= x"00ce5b04";
		wait for Clk_period;
		Addr <=  "00000110000010";
		Trees_din <= x"ff8c062d";
		wait for Clk_period;
		Addr <=  "00000110000011";
		Trees_din <= x"02fa4c04";
		wait for Clk_period;
		Addr <=  "00000110000100";
		Trees_din <= x"ffcd062d";
		wait for Clk_period;
		Addr <=  "00000110000101";
		Trees_din <= x"060d1804";
		wait for Clk_period;
		Addr <=  "00000110000110";
		Trees_din <= x"0021062d";
		wait for Clk_period;
		Addr <=  "00000110000111";
		Trees_din <= x"007d062d";
		wait for Clk_period;
		Addr <=  "00000110001000";
		Trees_din <= x"0123d704";
		wait for Clk_period;
		Addr <=  "00000110001001";
		Trees_din <= x"0091062d";
		wait for Clk_period;
		Addr <=  "00000110001010";
		Trees_din <= x"fff9062d";
		wait for Clk_period;
		Addr <=  "00000110001011";
		Trees_din <= x"060e1c14";
		wait for Clk_period;
		Addr <=  "00000110001100";
		Trees_din <= x"06047104";
		wait for Clk_period;
		Addr <=  "00000110001101";
		Trees_din <= x"ff690681";
		wait for Clk_period;
		Addr <=  "00000110001110";
		Trees_din <= x"00f45908";
		wait for Clk_period;
		Addr <=  "00000110001111";
		Trees_din <= x"0201bc04";
		wait for Clk_period;
		Addr <=  "00000110010000";
		Trees_din <= x"fffa0681";
		wait for Clk_period;
		Addr <=  "00000110010001";
		Trees_din <= x"ff840681";
		wait for Clk_period;
		Addr <=  "00000110010010";
		Trees_din <= x"04018604";
		wait for Clk_period;
		Addr <=  "00000110010011";
		Trees_din <= x"006e0681";
		wait for Clk_period;
		Addr <=  "00000110010100";
		Trees_din <= x"ffd90681";
		wait for Clk_period;
		Addr <=  "00000110010101";
		Trees_din <= x"02145114";
		wait for Clk_period;
		Addr <=  "00000110010110";
		Trees_din <= x"011cba0c";
		wait for Clk_period;
		Addr <=  "00000110010111";
		Trees_din <= x"07005b04";
		wait for Clk_period;
		Addr <=  "00000110011000";
		Trees_din <= x"00930681";
		wait for Clk_period;
		Addr <=  "00000110011001";
		Trees_din <= x"05ffb204";
		wait for Clk_period;
		Addr <=  "00000110011010";
		Trees_din <= x"00670681";
		wait for Clk_period;
		Addr <=  "00000110011011";
		Trees_din <= x"ffe60681";
		wait for Clk_period;
		Addr <=  "00000110011100";
		Trees_din <= x"1c004004";
		wait for Clk_period;
		Addr <=  "00000110011101";
		Trees_din <= x"ffe20681";
		wait for Clk_period;
		Addr <=  "00000110011110";
		Trees_din <= x"003c0681";
		wait for Clk_period;
		Addr <=  "00000110011111";
		Trees_din <= x"ffe20681";
		wait for Clk_period;
		Addr <=  "00000110100000";
		Trees_din <= x"0609350c";
		wait for Clk_period;
		Addr <=  "00000110100001";
		Trees_din <= x"11000004";
		wait for Clk_period;
		Addr <=  "00000110100010";
		Trees_din <= x"001006cd";
		wait for Clk_period;
		Addr <=  "00000110100011";
		Trees_din <= x"06080304";
		wait for Clk_period;
		Addr <=  "00000110100100";
		Trees_din <= x"ff6a06cd";
		wait for Clk_period;
		Addr <=  "00000110100101";
		Trees_din <= x"ffeb06cd";
		wait for Clk_period;
		Addr <=  "00000110100110";
		Trees_din <= x"060f950c";
		wait for Clk_period;
		Addr <=  "00000110100111";
		Trees_din <= x"04040104";
		wait for Clk_period;
		Addr <=  "00000110101000";
		Trees_din <= x"004806cd";
		wait for Clk_period;
		Addr <=  "00000110101001";
		Trees_din <= x"05feb204";
		wait for Clk_period;
		Addr <=  "00000110101010";
		Trees_din <= x"000306cd";
		wait for Clk_period;
		Addr <=  "00000110101011";
		Trees_din <= x"ff9706cd";
		wait for Clk_period;
		Addr <=  "00000110101100";
		Trees_din <= x"0123d70c";
		wait for Clk_period;
		Addr <=  "00000110101101";
		Trees_din <= x"07005b04";
		wait for Clk_period;
		Addr <=  "00000110101110";
		Trees_din <= x"008b06cd";
		wait for Clk_period;
		Addr <=  "00000110101111";
		Trees_din <= x"05fdc404";
		wait for Clk_period;
		Addr <=  "00000110110000";
		Trees_din <= x"005f06cd";
		wait for Clk_period;
		Addr <=  "00000110110001";
		Trees_din <= x"ffdd06cd";
		wait for Clk_period;
		Addr <=  "00000110110010";
		Trees_din <= x"ffee06cd";
		wait for Clk_period;
		Addr <=  "00000110110011";
		Trees_din <= x"060e1c14";
		wait for Clk_period;
		Addr <=  "00000110110100";
		Trees_din <= x"06047104";
		wait for Clk_period;
		Addr <=  "00000110110101";
		Trees_din <= x"ff6c0719";
		wait for Clk_period;
		Addr <=  "00000110110110";
		Trees_din <= x"00f45908";
		wait for Clk_period;
		Addr <=  "00000110110111";
		Trees_din <= x"0201bc04";
		wait for Clk_period;
		Addr <=  "00000110111000";
		Trees_din <= x"fff80719";
		wait for Clk_period;
		Addr <=  "00000110111001";
		Trees_din <= x"ff900719";
		wait for Clk_period;
		Addr <=  "00000110111010";
		Trees_din <= x"03fea104";
		wait for Clk_period;
		Addr <=  "00000110111011";
		Trees_din <= x"00630719";
		wait for Clk_period;
		Addr <=  "00000110111100";
		Trees_din <= x"ffea0719";
		wait for Clk_period;
		Addr <=  "00000110111101";
		Trees_din <= x"02145110";
		wait for Clk_period;
		Addr <=  "00000110111110";
		Trees_din <= x"011cba0c";
		wait for Clk_period;
		Addr <=  "00000110111111";
		Trees_din <= x"07005b04";
		wait for Clk_period;
		Addr <=  "00000111000000";
		Trees_din <= x"008d0719";
		wait for Clk_period;
		Addr <=  "00000111000001";
		Trees_din <= x"05ffb204";
		wait for Clk_period;
		Addr <=  "00000111000010";
		Trees_din <= x"00580719";
		wait for Clk_period;
		Addr <=  "00000111000011";
		Trees_din <= x"ffec0719";
		wait for Clk_period;
		Addr <=  "00000111000100";
		Trees_din <= x"00150719";
		wait for Clk_period;
		Addr <=  "00000111000101";
		Trees_din <= x"ffe70719";
		wait for Clk_period;
		Addr <=  "00000111000110";
		Trees_din <= x"060e1c14";
		wait for Clk_period;
		Addr <=  "00000111000111";
		Trees_din <= x"06047104";
		wait for Clk_period;
		Addr <=  "00000111001000";
		Trees_din <= x"ff6d0765";
		wait for Clk_period;
		Addr <=  "00000111001001";
		Trees_din <= x"0403c808";
		wait for Clk_period;
		Addr <=  "00000111001010";
		Trees_din <= x"0a01c204";
		wait for Clk_period;
		Addr <=  "00000111001011";
		Trees_din <= x"fff70765";
		wait for Clk_period;
		Addr <=  "00000111001100";
		Trees_din <= x"004d0765";
		wait for Clk_period;
		Addr <=  "00000111001101";
		Trees_din <= x"0f015604";
		wait for Clk_period;
		Addr <=  "00000111001110";
		Trees_din <= x"ffee0765";
		wait for Clk_period;
		Addr <=  "00000111001111";
		Trees_din <= x"ff940765";
		wait for Clk_period;
		Addr <=  "00000111010000";
		Trees_din <= x"02145110";
		wait for Clk_period;
		Addr <=  "00000111010001";
		Trees_din <= x"011cba0c";
		wait for Clk_period;
		Addr <=  "00000111010010";
		Trees_din <= x"07005b04";
		wait for Clk_period;
		Addr <=  "00000111010011";
		Trees_din <= x"00890765";
		wait for Clk_period;
		Addr <=  "00000111010100";
		Trees_din <= x"13fc8304";
		wait for Clk_period;
		Addr <=  "00000111010101";
		Trees_din <= x"fffa0765";
		wait for Clk_period;
		Addr <=  "00000111010110";
		Trees_din <= x"00490765";
		wait for Clk_period;
		Addr <=  "00000111010111";
		Trees_din <= x"00130765";
		wait for Clk_period;
		Addr <=  "00000111011000";
		Trees_din <= x"ffec0765";
		wait for Clk_period;
		Addr <=  "00000111011001";
		Trees_din <= x"060f9514";
		wait for Clk_period;
		Addr <=  "00000111011010";
		Trees_din <= x"06047104";
		wait for Clk_period;
		Addr <=  "00000111011011";
		Trees_din <= x"ff6f07a9";
		wait for Clk_period;
		Addr <=  "00000111011100";
		Trees_din <= x"04040108";
		wait for Clk_period;
		Addr <=  "00000111011101";
		Trees_din <= x"1a003e04";
		wait for Clk_period;
		Addr <=  "00000111011110";
		Trees_din <= x"004c07a9";
		wait for Clk_period;
		Addr <=  "00000111011111";
		Trees_din <= x"fffe07a9";
		wait for Clk_period;
		Addr <=  "00000111100000";
		Trees_din <= x"05feb204";
		wait for Clk_period;
		Addr <=  "00000111100001";
		Trees_din <= x"ffef07a9";
		wait for Clk_period;
		Addr <=  "00000111100010";
		Trees_din <= x"ff9a07a9";
		wait for Clk_period;
		Addr <=  "00000111100011";
		Trees_din <= x"011fa00c";
		wait for Clk_period;
		Addr <=  "00000111100100";
		Trees_din <= x"07005b04";
		wait for Clk_period;
		Addr <=  "00000111100101";
		Trees_din <= x"008207a9";
		wait for Clk_period;
		Addr <=  "00000111100110";
		Trees_din <= x"0d020f04";
		wait for Clk_period;
		Addr <=  "00000111100111";
		Trees_din <= x"003407a9";
		wait for Clk_period;
		Addr <=  "00000111101000";
		Trees_din <= x"fff307a9";
		wait for Clk_period;
		Addr <=  "00000111101001";
		Trees_din <= x"fffc07a9";
		wait for Clk_period;
		Addr <=  "00000111101010";
		Trees_din <= x"0609350c";
		wait for Clk_period;
		Addr <=  "00000111101011";
		Trees_din <= x"06047104";
		wait for Clk_period;
		Addr <=  "00000111101100";
		Trees_din <= x"ff7207e5";
		wait for Clk_period;
		Addr <=  "00000111101101";
		Trees_din <= x"01feba04";
		wait for Clk_period;
		Addr <=  "00000111101110";
		Trees_din <= x"002a07e5";
		wait for Clk_period;
		Addr <=  "00000111101111";
		Trees_din <= x"ffaf07e5";
		wait for Clk_period;
		Addr <=  "00000111110000";
		Trees_din <= x"0613800c";
		wait for Clk_period;
		Addr <=  "00000111110001";
		Trees_din <= x"00d71804";
		wait for Clk_period;
		Addr <=  "00000111110010";
		Trees_din <= x"ffab07e5";
		wait for Clk_period;
		Addr <=  "00000111110011";
		Trees_din <= x"0f027804";
		wait for Clk_period;
		Addr <=  "00000111110100";
		Trees_din <= x"005007e5";
		wait for Clk_period;
		Addr <=  "00000111110101";
		Trees_din <= x"fff007e5";
		wait for Clk_period;
		Addr <=  "00000111110110";
		Trees_din <= x"0413db04";
		wait for Clk_period;
		Addr <=  "00000111110111";
		Trees_din <= x"007807e5";
		wait for Clk_period;
		Addr <=  "00000111111000";
		Trees_din <= x"002007e5";
		wait for Clk_period;
		Addr <=  "00000111111001";
		Trees_din <= x"060f9514";
		wait for Clk_period;
		Addr <=  "00000111111010";
		Trees_din <= x"06047104";
		wait for Clk_period;
		Addr <=  "00000111111011";
		Trees_din <= x"ff750821";
		wait for Clk_period;
		Addr <=  "00000111111100";
		Trees_din <= x"04040108";
		wait for Clk_period;
		Addr <=  "00000111111101";
		Trees_din <= x"03fe5704";
		wait for Clk_period;
		Addr <=  "00000111111110";
		Trees_din <= x"003c0821";
		wait for Clk_period;
		Addr <=  "00000111111111";
		Trees_din <= x"fff90821";
		wait for Clk_period;
		Addr <=  "00001000000000";
		Trees_din <= x"05feb204";
		wait for Clk_period;
		Addr <=  "00001000000001";
		Trees_din <= x"ffed0821";
		wait for Clk_period;
		Addr <=  "00001000000010";
		Trees_din <= x"ffa70821";
		wait for Clk_period;
		Addr <=  "00001000000011";
		Trees_din <= x"0413db08";
		wait for Clk_period;
		Addr <=  "00001000000100";
		Trees_din <= x"07005b04";
		wait for Clk_period;
		Addr <=  "00001000000101";
		Trees_din <= x"00730821";
		wait for Clk_period;
		Addr <=  "00001000000110";
		Trees_din <= x"00120821";
		wait for Clk_period;
		Addr <=  "00001000000111";
		Trees_din <= x"00070821";
		wait for Clk_period;
		Addr <=  "00001000001000";
		Trees_din <= x"06093508";
		wait for Clk_period;
		Addr <=  "00001000001001";
		Trees_din <= x"06047104";
		wait for Clk_period;
		Addr <=  "00001000001010";
		Trees_din <= x"ff78084d";
		wait for Clk_period;
		Addr <=  "00001000001011";
		Trees_din <= x"ffe5084d";
		wait for Clk_period;
		Addr <=  "00001000001100";
		Trees_din <= x"0614d40c";
		wait for Clk_period;
		Addr <=  "00001000001101";
		Trees_din <= x"00d25d04";
		wait for Clk_period;
		Addr <=  "00001000001110";
		Trees_din <= x"ffb0084d";
		wait for Clk_period;
		Addr <=  "00001000001111";
		Trees_din <= x"05ff3a04";
		wait for Clk_period;
		Addr <=  "00001000010000";
		Trees_din <= x"0048084d";
		wait for Clk_period;
		Addr <=  "00001000010001";
		Trees_din <= x"fff5084d";
		wait for Clk_period;
		Addr <=  "00001000010010";
		Trees_din <= x"0068084d";
		wait for Clk_period;
		Addr <=  "00001000010011";
		Trees_din <= x"060e1c10";
		wait for Clk_period;
		Addr <=  "00001000010100";
		Trees_din <= x"06047104";
		wait for Clk_period;
		Addr <=  "00001000010101";
		Trees_din <= x"ff7c0881";
		wait for Clk_period;
		Addr <=  "00001000010110";
		Trees_din <= x"18003104";
		wait for Clk_period;
		Addr <=  "00001000010111";
		Trees_din <= x"00300881";
		wait for Clk_period;
		Addr <=  "00001000011000";
		Trees_din <= x"00f45904";
		wait for Clk_period;
		Addr <=  "00001000011001";
		Trees_din <= x"ffae0881";
		wait for Clk_period;
		Addr <=  "00001000011010";
		Trees_din <= x"fff90881";
		wait for Clk_period;
		Addr <=  "00001000011011";
		Trees_din <= x"061cb508";
		wait for Clk_period;
		Addr <=  "00001000011100";
		Trees_din <= x"00c00004";
		wait for Clk_period;
		Addr <=  "00001000011101";
		Trees_din <= x"ffb60881";
		wait for Clk_period;
		Addr <=  "00001000011110";
		Trees_din <= x"00580881";
		wait for Clk_period;
		Addr <=  "00001000011111";
		Trees_din <= x"00760881";
		wait for Clk_period;
		Addr <=  "00001000100000";
		Trees_din <= x"060f950c";
		wait for Clk_period;
		Addr <=  "00001000100001";
		Trees_din <= x"06047104";
		wait for Clk_period;
		Addr <=  "00001000100010";
		Trees_din <= x"ff8008ad";
		wait for Clk_period;
		Addr <=  "00001000100011";
		Trees_din <= x"04040104";
		wait for Clk_period;
		Addr <=  "00001000100100";
		Trees_din <= x"001e08ad";
		wait for Clk_period;
		Addr <=  "00001000100101";
		Trees_din <= x"ffbe08ad";
		wait for Clk_period;
		Addr <=  "00001000100110";
		Trees_din <= x"061cb508";
		wait for Clk_period;
		Addr <=  "00001000100111";
		Trees_din <= x"00c00004";
		wait for Clk_period;
		Addr <=  "00001000101000";
		Trees_din <= x"ffbf08ad";
		wait for Clk_period;
		Addr <=  "00001000101001";
		Trees_din <= x"005408ad";
		wait for Clk_period;
		Addr <=  "00001000101010";
		Trees_din <= x"007108ad";
		wait for Clk_period;
		Addr <=  "00001000101011";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00001000101100";
		Trees_din <= x"060e1c0c";
		wait for Clk_period;
		Addr <=  "00001000101101";
		Trees_din <= x"06047104";
		wait for Clk_period;
		Addr <=  "00001000101110";
		Trees_din <= x"ff8508dd";
		wait for Clk_period;
		Addr <=  "00001000101111";
		Trees_din <= x"00f45904";
		wait for Clk_period;
		Addr <=  "00001000110000";
		Trees_din <= x"ffc208dd";
		wait for Clk_period;
		Addr <=  "00001000110001";
		Trees_din <= x"001a08dd";
		wait for Clk_period;
		Addr <=  "00001000110010";
		Trees_din <= x"0614d404";
		wait for Clk_period;
		Addr <=  "00001000110011";
		Trees_din <= x"000508dd";
		wait for Clk_period;
		Addr <=  "00001000110100";
		Trees_din <= x"061cb504";
		wait for Clk_period;
		Addr <=  "00001000110101";
		Trees_din <= x"002508dd";
		wait for Clk_period;
		Addr <=  "00001000110110";
		Trees_din <= x"006c08dd";
		wait for Clk_period;
		Addr <=  "00001000110111";
		Trees_din <= x"060f950c";
		wait for Clk_period;
		Addr <=  "00001000111000";
		Trees_din <= x"06047104";
		wait for Clk_period;
		Addr <=  "00001000111001";
		Trees_din <= x"ff8a0901";
		wait for Clk_period;
		Addr <=  "00001000111010";
		Trees_din <= x"0a02ce04";
		wait for Clk_period;
		Addr <=  "00001000111011";
		Trees_din <= x"ffc90901";
		wait for Clk_period;
		Addr <=  "00001000111100";
		Trees_din <= x"00220901";
		wait for Clk_period;
		Addr <=  "00001000111101";
		Trees_din <= x"07005b04";
		wait for Clk_period;
		Addr <=  "00001000111110";
		Trees_din <= x"00550901";
		wait for Clk_period;
		Addr <=  "00001000111111";
		Trees_din <= x"00010901";
		wait for Clk_period;
		Addr <=  "00001001000000";
		Trees_din <= x"06138010";
		wait for Clk_period;
		Addr <=  "00001001000001";
		Trees_din <= x"06047104";
		wait for Clk_period;
		Addr <=  "00001001000010";
		Trees_din <= x"ff8f092d";
		wait for Clk_period;
		Addr <=  "00001001000011";
		Trees_din <= x"0207cc08";
		wait for Clk_period;
		Addr <=  "00001001000100";
		Trees_din <= x"02ffbf04";
		wait for Clk_period;
		Addr <=  "00001001000101";
		Trees_din <= x"ffed092d";
		wait for Clk_period;
		Addr <=  "00001001000110";
		Trees_din <= x"002d092d";
		wait for Clk_period;
		Addr <=  "00001001000111";
		Trees_din <= x"ffb6092d";
		wait for Clk_period;
		Addr <=  "00001001001000";
		Trees_din <= x"061cb504";
		wait for Clk_period;
		Addr <=  "00001001001001";
		Trees_din <= x"001e092d";
		wait for Clk_period;
		Addr <=  "00001001001010";
		Trees_din <= x"0064092d";
		wait for Clk_period;
		Addr <=  "00001001001011";
		Trees_din <= x"060e1c08";
		wait for Clk_period;
		Addr <=  "00001001001100";
		Trees_din <= x"18003104";
		wait for Clk_period;
		Addr <=  "00001001001101";
		Trees_din <= x"fffd0951";
		wait for Clk_period;
		Addr <=  "00001001001110";
		Trees_din <= x"ffa20951";
		wait for Clk_period;
		Addr <=  "00001001001111";
		Trees_din <= x"061cb508";
		wait for Clk_period;
		Addr <=  "00001001010000";
		Trees_din <= x"00c02704";
		wait for Clk_period;
		Addr <=  "00001001010001";
		Trees_din <= x"ffc60951";
		wait for Clk_period;
		Addr <=  "00001001010010";
		Trees_din <= x"00480951";
		wait for Clk_period;
		Addr <=  "00001001010011";
		Trees_din <= x"00600951";
		wait for Clk_period;
		Addr <=  "00001001010100";
		Trees_din <= x"06093508";
		wait for Clk_period;
		Addr <=  "00001001010101";
		Trees_din <= x"06047104";
		wait for Clk_period;
		Addr <=  "00001001010110";
		Trees_din <= x"ff990975";
		wait for Clk_period;
		Addr <=  "00001001010111";
		Trees_din <= x"ffeb0975";
		wait for Clk_period;
		Addr <=  "00001001011000";
		Trees_din <= x"0615fc08";
		wait for Clk_period;
		Addr <=  "00001001011001";
		Trees_din <= x"05feb204";
		wait for Clk_period;
		Addr <=  "00001001011010";
		Trees_din <= x"00310975";
		wait for Clk_period;
		Addr <=  "00001001011011";
		Trees_din <= x"ffcd0975";
		wait for Clk_period;
		Addr <=  "00001001011100";
		Trees_din <= x"00500975";
		wait for Clk_period;
		Addr <=  "00001001011101";
		Trees_din <= x"060d1808";
		wait for Clk_period;
		Addr <=  "00001001011110";
		Trees_din <= x"1a003e04";
		wait for Clk_period;
		Addr <=  "00001001011111";
		Trees_din <= x"fff90999";
		wait for Clk_period;
		Addr <=  "00001001100000";
		Trees_din <= x"ffa40999";
		wait for Clk_period;
		Addr <=  "00001001100001";
		Trees_din <= x"05fe0104";
		wait for Clk_period;
		Addr <=  "00001001100010";
		Trees_din <= x"00570999";
		wait for Clk_period;
		Addr <=  "00001001100011";
		Trees_din <= x"13fcd204";
		wait for Clk_period;
		Addr <=  "00001001100100";
		Trees_din <= x"ffe60999";
		wait for Clk_period;
		Addr <=  "00001001100101";
		Trees_din <= x"00270999";
		wait for Clk_period;
		Addr <=  "00001001100110";
		Trees_din <= x"0613800c";
		wait for Clk_period;
		Addr <=  "00001001100111";
		Trees_din <= x"06047104";
		wait for Clk_period;
		Addr <=  "00001001101000";
		Trees_din <= x"ffa209bd";
		wait for Clk_period;
		Addr <=  "00001001101001";
		Trees_din <= x"02051104";
		wait for Clk_period;
		Addr <=  "00001001101010";
		Trees_din <= x"001809bd";
		wait for Clk_period;
		Addr <=  "00001001101011";
		Trees_din <= x"ffc909bd";
		wait for Clk_period;
		Addr <=  "00001001101100";
		Trees_din <= x"061cb504";
		wait for Clk_period;
		Addr <=  "00001001101101";
		Trees_din <= x"001609bd";
		wait for Clk_period;
		Addr <=  "00001001101110";
		Trees_din <= x"005709bd";
		wait for Clk_period;
		Addr <=  "00001001101111";
		Trees_din <= x"0613800c";
		wait for Clk_period;
		Addr <=  "00001001110000";
		Trees_din <= x"06047104";
		wait for Clk_period;
		Addr <=  "00001001110001";
		Trees_din <= x"ffa709e1";
		wait for Clk_period;
		Addr <=  "00001001110010";
		Trees_din <= x"04044704";
		wait for Clk_period;
		Addr <=  "00001001110011";
		Trees_din <= x"001c09e1";
		wait for Clk_period;
		Addr <=  "00001001110100";
		Trees_din <= x"ffd809e1";
		wait for Clk_period;
		Addr <=  "00001001110101";
		Trees_din <= x"061cb504";
		wait for Clk_period;
		Addr <=  "00001001110110";
		Trees_din <= x"001609e1";
		wait for Clk_period;
		Addr <=  "00001001110111";
		Trees_din <= x"005309e1";
		wait for Clk_period;
		Addr <=  "00001001111000";
		Trees_din <= x"060e1c08";
		wait for Clk_period;
		Addr <=  "00001001111001";
		Trees_din <= x"0a02ce04";
		wait for Clk_period;
		Addr <=  "00001001111010";
		Trees_din <= x"ffb309fd";
		wait for Clk_period;
		Addr <=  "00001001111011";
		Trees_din <= x"000009fd";
		wait for Clk_period;
		Addr <=  "00001001111100";
		Trees_din <= x"0615fc04";
		wait for Clk_period;
		Addr <=  "00001001111101";
		Trees_din <= x"000609fd";
		wait for Clk_period;
		Addr <=  "00001001111110";
		Trees_din <= x"004609fd";
		wait for Clk_period;
		Addr <=  "00001001111111";
		Trees_din <= x"06093504";
		wait for Clk_period;
		Addr <=  "00001010000000";
		Trees_din <= x"ffbc0a19";
		wait for Clk_period;
		Addr <=  "00001010000001";
		Trees_din <= x"05fe0104";
		wait for Clk_period;
		Addr <=  "00001010000010";
		Trees_din <= x"00450a19";
		wait for Clk_period;
		Addr <=  "00001010000011";
		Trees_din <= x"13fd0204";
		wait for Clk_period;
		Addr <=  "00001010000100";
		Trees_din <= x"ffeb0a19";
		wait for Clk_period;
		Addr <=  "00001010000101";
		Trees_din <= x"001d0a19";
		wait for Clk_period;
		Addr <=  "00001010000110";
		Trees_din <= x"0613800c";
		wait for Clk_period;
		Addr <=  "00001010000111";
		Trees_din <= x"06047104";
		wait for Clk_period;
		Addr <=  "00001010001000";
		Trees_din <= x"ffb30a35";
		wait for Clk_period;
		Addr <=  "00001010001001";
		Trees_din <= x"04044704";
		wait for Clk_period;
		Addr <=  "00001010001010";
		Trees_din <= x"001c0a35";
		wait for Clk_period;
		Addr <=  "00001010001011";
		Trees_din <= x"ffdd0a35";
		wait for Clk_period;
		Addr <=  "00001010001100";
		Trees_din <= x"003d0a35";
		wait for Clk_period;
		Addr <=  "00001010001101";
		Trees_din <= x"060e1c08";
		wait for Clk_period;
		Addr <=  "00001010001110";
		Trees_din <= x"1d00db04";
		wait for Clk_period;
		Addr <=  "00001010001111";
		Trees_din <= x"ffbf0a51";
		wait for Clk_period;
		Addr <=  "00001010010000";
		Trees_din <= x"fffc0a51";
		wait for Clk_period;
		Addr <=  "00001010010001";
		Trees_din <= x"11021d04";
		wait for Clk_period;
		Addr <=  "00001010010010";
		Trees_din <= x"00400a51";
		wait for Clk_period;
		Addr <=  "00001010010011";
		Trees_din <= x"00040a51";
		wait for Clk_period;
		Addr <=  "00001010010100";
		Trees_din <= x"0614d40c";
		wait for Clk_period;
		Addr <=  "00001010010101";
		Trees_din <= x"0501ea08";
		wait for Clk_period;
		Addr <=  "00001010010110";
		Trees_din <= x"1b01aa04";
		wait for Clk_period;
		Addr <=  "00001010010111";
		Trees_din <= x"00180a6d";
		wait for Clk_period;
		Addr <=  "00001010011000";
		Trees_din <= x"ffe40a6d";
		wait for Clk_period;
		Addr <=  "00001010011001";
		Trees_din <= x"ffbb0a6d";
		wait for Clk_period;
		Addr <=  "00001010011010";
		Trees_din <= x"003a0a6d";
		wait for Clk_period;
		Addr <=  "00001010011011";
		Trees_din <= x"060af004";
		wait for Clk_period;
		Addr <=  "00001010011100";
		Trees_din <= x"ffca0a81";
		wait for Clk_period;
		Addr <=  "00001010011101";
		Trees_din <= x"05fe0104";
		wait for Clk_period;
		Addr <=  "00001010011110";
		Trees_din <= x"00410a81";
		wait for Clk_period;
		Addr <=  "00001010011111";
		Trees_din <= x"00030a81";
		wait for Clk_period;
		Addr <=  "00001010100000";
		Trees_din <= x"06080304";
		wait for Clk_period;
		Addr <=  "00001010100001";
		Trees_din <= x"ffc70a9d";
		wait for Clk_period;
		Addr <=  "00001010100010";
		Trees_din <= x"05fe0104";
		wait for Clk_period;
		Addr <=  "00001010100011";
		Trees_din <= x"00380a9d";
		wait for Clk_period;
		Addr <=  "00001010100100";
		Trees_din <= x"13fd0204";
		wait for Clk_period;
		Addr <=  "00001010100101";
		Trees_din <= x"ffed0a9d";
		wait for Clk_period;
		Addr <=  "00001010100110";
		Trees_din <= x"00190a9d";
		wait for Clk_period;
		Addr <=  "00001010100111";
		Trees_din <= x"0615fc08";
		wait for Clk_period;
		Addr <=  "00001010101000";
		Trees_din <= x"1400cd04";
		wait for Clk_period;
		Addr <=  "00001010101001";
		Trees_din <= x"000d0ab1";
		wait for Clk_period;
		Addr <=  "00001010101010";
		Trees_din <= x"ffd00ab1";
		wait for Clk_period;
		Addr <=  "00001010101011";
		Trees_din <= x"00390ab1";
		wait for Clk_period;
		Addr <=  "00001010101100";
		Trees_din <= x"060e1c04";
		wait for Clk_period;
		Addr <=  "00001010101101";
		Trees_din <= x"ffd90ac5";
		wait for Clk_period;
		Addr <=  "00001010101110";
		Trees_din <= x"1101ce04";
		wait for Clk_period;
		Addr <=  "00001010101111";
		Trees_din <= x"00380ac5";
		wait for Clk_period;
		Addr <=  "00001010110000";
		Trees_din <= x"00040ac5";
		wait for Clk_period;
		Addr <=  "00001010110001";
		Trees_din <= x"0a029908";
		wait for Clk_period;
		Addr <=  "00001010110010";
		Trees_din <= x"060f9504";
		wait for Clk_period;
		Addr <=  "00001010110011";
		Trees_din <= x"ffcb0ad9";
		wait for Clk_period;
		Addr <=  "00001010110100";
		Trees_din <= x"00150ad9";
		wait for Clk_period;
		Addr <=  "00001010110101";
		Trees_din <= x"00230ad9";
		wait for Clk_period;
		Addr <=  "00001010110110";
		Trees_din <= x"0a029908";
		wait for Clk_period;
		Addr <=  "00001010110111";
		Trees_din <= x"060e1c04";
		wait for Clk_period;
		Addr <=  "00001010111000";
		Trees_din <= x"ffcd0aed";
		wait for Clk_period;
		Addr <=  "00001010111001";
		Trees_din <= x"00130aed";
		wait for Clk_period;
		Addr <=  "00001010111010";
		Trees_din <= x"00200aed";
		wait for Clk_period;
		Addr <=  "00001010111011";
		Trees_din <= x"05fde404";
		wait for Clk_period;
		Addr <=  "00001010111100";
		Trees_din <= x"00210b01";
		wait for Clk_period;
		Addr <=  "00001010111101";
		Trees_din <= x"0b003d04";
		wait for Clk_period;
		Addr <=  "00001010111110";
		Trees_din <= x"00140b01";
		wait for Clk_period;
		Addr <=  "00001010111111";
		Trees_din <= x"ffd80b01";
		wait for Clk_period;
		Addr <=  "00001011000000";
		Trees_din <= x"0615fc08";
		wait for Clk_period;
		Addr <=  "00001011000001";
		Trees_din <= x"05feb204";
		wait for Clk_period;
		Addr <=  "00001011000010";
		Trees_din <= x"00080b15";
		wait for Clk_period;
		Addr <=  "00001011000011";
		Trees_din <= x"ffd40b15";
		wait for Clk_period;
		Addr <=  "00001011000100";
		Trees_din <= x"00340b15";
		wait for Clk_period;
		Addr <=  "00001011000101";
		Trees_din <= x"17003d04";
		wait for Clk_period;
		Addr <=  "00001011000110";
		Trees_din <= x"001f0b29";
		wait for Clk_period;
		Addr <=  "00001011000111";
		Trees_din <= x"11020904";
		wait for Clk_period;
		Addr <=  "00001011001000";
		Trees_din <= x"00080b29";
		wait for Clk_period;
		Addr <=  "00001011001001";
		Trees_din <= x"ffe00b29";
		wait for Clk_period;
		Addr <=  "00001011001010";
		Trees_din <= x"060e1c04";
		wait for Clk_period;
		Addr <=  "00001011001011";
		Trees_din <= x"ffdc0b35";
		wait for Clk_period;
		Addr <=  "00001011001100";
		Trees_din <= x"00260b35";
		wait for Clk_period;
		Addr <=  "00001011001101";
		Trees_din <= x"0a029908";
		wait for Clk_period;
		Addr <=  "00001011001110";
		Trees_din <= x"14030b04";
		wait for Clk_period;
		Addr <=  "00001011001111";
		Trees_din <= x"ffe50b49";
		wait for Clk_period;
		Addr <=  "00001011010000";
		Trees_din <= x"00020b49";
		wait for Clk_period;
		Addr <=  "00001011010001";
		Trees_din <= x"001b0b49";
		wait for Clk_period;
		Addr <=  "00001011010010";
		Trees_din <= x"05fde404";
		wait for Clk_period;
		Addr <=  "00001011010011";
		Trees_din <= x"001c0b5d";
		wait for Clk_period;
		Addr <=  "00001011010100";
		Trees_din <= x"0b003d04";
		wait for Clk_period;
		Addr <=  "00001011010101";
		Trees_din <= x"00110b5d";
		wait for Clk_period;
		Addr <=  "00001011010110";
		Trees_din <= x"ffdc0b5d";
		wait for Clk_period;
		Addr <=  "00001011010111";
		Trees_din <= x"0614d408";
		wait for Clk_period;
		Addr <=  "00001011011000";
		Trees_din <= x"05ff8704";
		wait for Clk_period;
		Addr <=  "00001011011001";
		Trees_din <= x"00010b71";
		wait for Clk_period;
		Addr <=  "00001011011010";
		Trees_din <= x"ffd50b71";
		wait for Clk_period;
		Addr <=  "00001011011011";
		Trees_din <= x"002f0b71";
		wait for Clk_period;
		Addr <=  "00001011011100";
		Trees_din <= x"17003d04";
		wait for Clk_period;
		Addr <=  "00001011011101";
		Trees_din <= x"001b0b85";
		wait for Clk_period;
		Addr <=  "00001011011110";
		Trees_din <= x"0eff7d04";
		wait for Clk_period;
		Addr <=  "00001011011111";
		Trees_din <= x"ffe20b85";
		wait for Clk_period;
		Addr <=  "00001011100000";
		Trees_din <= x"000a0b85";
		wait for Clk_period;
		Addr <=  "00001011100001";
		Trees_din <= x"17003d04";
		wait for Clk_period;
		Addr <=  "00001011100010";
		Trees_din <= x"00190b99";
		wait for Clk_period;
		Addr <=  "00001011100011";
		Trees_din <= x"0eff7d04";
		wait for Clk_period;
		Addr <=  "00001011100100";
		Trees_din <= x"ffe50b99";
		wait for Clk_period;
		Addr <=  "00001011100101";
		Trees_din <= x"00090b99";
		wait for Clk_period;
		Addr <=  "00001011100110";
		Trees_din <= x"060af004";
		wait for Clk_period;
		Addr <=  "00001011100111";
		Trees_din <= x"ffd50bad";
		wait for Clk_period;
		Addr <=  "00001011101000";
		Trees_din <= x"13fd0204";
		wait for Clk_period;
		Addr <=  "00001011101001";
		Trees_din <= x"00050bad";
		wait for Clk_period;
		Addr <=  "00001011101010";
		Trees_din <= x"00290bad";
		wait for Clk_period;
		Addr <=  "00001011101011";
		Trees_din <= x"05fde404";
		wait for Clk_period;
		Addr <=  "00001011101100";
		Trees_din <= x"001a0bc1";
		wait for Clk_period;
		Addr <=  "00001011101101";
		Trees_din <= x"0b003904";
		wait for Clk_period;
		Addr <=  "00001011101110";
		Trees_din <= x"000e0bc1";
		wait for Clk_period;
		Addr <=  "00001011101111";
		Trees_din <= x"ffdf0bc1";
		wait for Clk_period;
		Addr <=  "00001011110000";
		Trees_din <= x"05fde404";
		wait for Clk_period;
		Addr <=  "00001011110001";
		Trees_din <= x"00180bd5";
		wait for Clk_period;
		Addr <=  "00001011110010";
		Trees_din <= x"0b003904";
		wait for Clk_period;
		Addr <=  "00001011110011";
		Trees_din <= x"000c0bd5";
		wait for Clk_period;
		Addr <=  "00001011110100";
		Trees_din <= x"ffe20bd5";
		wait for Clk_period;
		Addr <=  "00001011110101";
		Trees_din <= x"060e1c04";
		wait for Clk_period;
		Addr <=  "00001011110110";
		Trees_din <= x"ffdc0be1";
		wait for Clk_period;
		Addr <=  "00001011110111";
		Trees_din <= x"00230be1";
		wait for Clk_period;
		Addr <=  "00001011111000";
		Trees_din <= x"17003d04";
		wait for Clk_period;
		Addr <=  "00001011111001";
		Trees_din <= x"00160bf5";
		wait for Clk_period;
		Addr <=  "00001011111010";
		Trees_din <= x"0eff7d04";
		wait for Clk_period;
		Addr <=  "00001011111011";
		Trees_din <= x"ffe50bf5";
		wait for Clk_period;
		Addr <=  "00001011111100";
		Trees_din <= x"00090bf5";
		wait for Clk_period;
		Addr <=  "00001011111101";
		Trees_din <= x"05feb204";
		wait for Clk_period;
		Addr <=  "00001011111110";
		Trees_din <= x"00130c01";
		wait for Clk_period;
		Addr <=  "00001011111111";
		Trees_din <= x"fff30c01";
		wait for Clk_period;
		Addr <=  "00001100000000";
		Trees_din <= x"00f01304";
		wait for Clk_period;
		Addr <=  "00001100000001";
		Trees_din <= x"000f0c0d";
		wait for Clk_period;
		Addr <=  "00001100000010";
		Trees_din <= x"ffeb0c0d";
		wait for Clk_period;
		Addr <=  "00001100000011";
		Trees_din <= x"1b015104";
		wait for Clk_period;
		Addr <=  "00001100000100";
		Trees_din <= x"00120c19";
		wait for Clk_period;
		Addr <=  "00001100000101";
		Trees_din <= x"fff20c19";
		wait for Clk_period;
		Addr <=  "00001100000110";
		Trees_din <= x"0eff8c04";
		wait for Clk_period;
		Addr <=  "00001100000111";
		Trees_din <= x"fff10c25";
		wait for Clk_period;
		Addr <=  "00001100001000";
		Trees_din <= x"00110c25";
		wait for Clk_period;
		Addr <=  "00001100001001";
		Trees_din <= x"0a029904";
		wait for Clk_period;
		Addr <=  "00001100001010";
		Trees_din <= x"fff30c31";
		wait for Clk_period;
		Addr <=  "00001100001011";
		Trees_din <= x"00110c31";
		wait for Clk_period;
		Addr <=  "00001100001100";
		Trees_din <= x"06138004";
		wait for Clk_period;
		Addr <=  "00001100001101";
		Trees_din <= x"ffe30c3d";
		wait for Clk_period;
		Addr <=  "00001100001110";
		Trees_din <= x"00280c3d";
		wait for Clk_period;
		Addr <=  "00001100001111";
		Trees_din <= x"05feb204";
		wait for Clk_period;
		Addr <=  "00001100010000";
		Trees_din <= x"00120c49";
		wait for Clk_period;
		Addr <=  "00001100010001";
		Trees_din <= x"fff30c49";
		wait for Clk_period;
		Addr <=  "00001100010010";
		Trees_din <= x"19009b04";
		wait for Clk_period;
		Addr <=  "00001100010011";
		Trees_din <= x"fff40c55";
		wait for Clk_period;
		Addr <=  "00001100010100";
		Trees_din <= x"00110c55";
		wait for Clk_period;
		Addr <=  "00001100010101";
		Trees_din <= x"00e76404";
		wait for Clk_period;
		Addr <=  "00001100010110";
		Trees_din <= x"000e0c61";
		wait for Clk_period;
		Addr <=  "00001100010111";
		Trees_din <= x"fff00c61";
		wait for Clk_period;
		Addr <=  "00001100011000";
		Trees_din <= x"15028204";
		wait for Clk_period;
		Addr <=  "00001100011001";
		Trees_din <= x"000f0c6d";
		wait for Clk_period;
		Addr <=  "00001100011010";
		Trees_din <= x"fff20c6d";
		wait for Clk_period;
		Addr <=  "00001100011011";
		Trees_din <= x"05feb204";
		wait for Clk_period;
		Addr <=  "00001100011100";
		Trees_din <= x"00110c79";
		wait for Clk_period;
		Addr <=  "00001100011101";
		Trees_din <= x"fff40c79";
		wait for Clk_period;
		Addr <=  "00001100011110";
		Trees_din <= x"06138004";
		wait for Clk_period;
		Addr <=  "00001100011111";
		Trees_din <= x"ffe40c85";
		wait for Clk_period;
		Addr <=  "00001100100000";
		Trees_din <= x"00270c85";
		wait for Clk_period;
		Addr <=  "00001100100001";
		Trees_din <= x"1b015104";
		wait for Clk_period;
		Addr <=  "00001100100010";
		Trees_din <= x"00100c91";
		wait for Clk_period;
		Addr <=  "00001100100011";
		Trees_din <= x"fff40c91";
		wait for Clk_period;
		Addr <=  "00001100100100";
		Trees_din <= x"05feb204";
		wait for Clk_period;
		Addr <=  "00001100100101";
		Trees_din <= x"00100c9d";
		wait for Clk_period;
		Addr <=  "00001100100110";
		Trees_din <= x"fff50c9d";
		wait for Clk_period;
		Addr <=  "00001100100111";
		Trees_din <= x"00e76404";
		wait for Clk_period;
		Addr <=  "00001100101000";
		Trees_din <= x"000d0ca9";
		wait for Clk_period;
		Addr <=  "00001100101001";
		Trees_din <= x"fff20ca9";
		wait for Clk_period;
		Addr <=  "00001100101010";
		Trees_din <= x"19009d04";
		wait for Clk_period;
		Addr <=  "00001100101011";
		Trees_din <= x"fff40cb5";
		wait for Clk_period;
		Addr <=  "00001100101100";
		Trees_din <= x"00110cb5";
		wait for Clk_period;
		Addr <=  "00001100101101";
		Trees_din <= x"13027104";
		wait for Clk_period;
		Addr <=  "00001100101110";
		Trees_din <= x"fff50cc1";
		wait for Clk_period;
		Addr <=  "00001100101111";
		Trees_din <= x"00100cc1";
		wait for Clk_period;
		Addr <=  "00001100110000";
		Trees_din <= x"05feb204";
		wait for Clk_period;
		Addr <=  "00001100110001";
		Trees_din <= x"00100ccd";
		wait for Clk_period;
		Addr <=  "00001100110010";
		Trees_din <= x"fff50ccd";
		wait for Clk_period;
		Addr <=  "00001100110011";
		Trees_din <= x"0eff7d04";
		wait for Clk_period;
		Addr <=  "00001100110100";
		Trees_din <= x"fff40cd9";
		wait for Clk_period;
		Addr <=  "00001100110101";
		Trees_din <= x"000e0cd9";
		wait for Clk_period;
		Addr <=  "00001100110110";
		Trees_din <= x"00e76404";
		wait for Clk_period;
		Addr <=  "00001100110111";
		Trees_din <= x"000c0ce5";
		wait for Clk_period;
		Addr <=  "00001100111000";
		Trees_din <= x"fff20ce5";
		wait for Clk_period;
		Addr <=  "00001100111001";
		Trees_din <= x"18003604";
		wait for Clk_period;
		Addr <=  "00001100111010";
		Trees_din <= x"000f0cf1";
		wait for Clk_period;
		Addr <=  "00001100111011";
		Trees_din <= x"fff40cf1";
		wait for Clk_period;
		Addr <=  "00001100111100";
		Trees_din <= x"13027104";
		wait for Clk_period;
		Addr <=  "00001100111101";
		Trees_din <= x"fff50cfd";
		wait for Clk_period;
		Addr <=  "00001100111110";
		Trees_din <= x"000e0cfd";
		wait for Clk_period;
		Addr <=  "00001100111111";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  3
        -----------
		Addr <=  "00000000000000";
		Trees_din <= x"01152c2c";
		wait for Clk_period;
		Addr <=  "00000000000001";
		Trees_din <= x"010e9020";
		wait for Clk_period;
		Addr <=  "00000000000010";
		Trees_din <= x"0105d604";
		wait for Clk_period;
		Addr <=  "00000000000011";
		Trees_din <= x"ff4e007d";
		wait for Clk_period;
		Addr <=  "00000000000100";
		Trees_din <= x"00f88410";
		wait for Clk_period;
		Addr <=  "00000000000101";
		Trees_din <= x"00f56608";
		wait for Clk_period;
		Addr <=  "00000000000110";
		Trees_din <= x"00e76404";
		wait for Clk_period;
		Addr <=  "00000000000111";
		Trees_din <= x"ff4f007d";
		wait for Clk_period;
		Addr <=  "00000000001000";
		Trees_din <= x"ffaa007d";
		wait for Clk_period;
		Addr <=  "00000000001001";
		Trees_din <= x"01081b04";
		wait for Clk_period;
		Addr <=  "00000000001010";
		Trees_din <= x"ff78007d";
		wait for Clk_period;
		Addr <=  "00000000001011";
		Trees_din <= x"0190007d";
		wait for Clk_period;
		Addr <=  "00000000001100";
		Trees_din <= x"020a6908";
		wait for Clk_period;
		Addr <=  "00000000001101";
		Trees_din <= x"0c014004";
		wait for Clk_period;
		Addr <=  "00000000001110";
		Trees_din <= x"031a007d";
		wait for Clk_period;
		Addr <=  "00000000001111";
		Trees_din <= x"010b007d";
		wait for Clk_period;
		Addr <=  "00000000010000";
		Trees_din <= x"ff85007d";
		wait for Clk_period;
		Addr <=  "00000000010001";
		Trees_din <= x"00dc8808";
		wait for Clk_period;
		Addr <=  "00000000010010";
		Trees_din <= x"00d71804";
		wait for Clk_period;
		Addr <=  "00000000010011";
		Trees_din <= x"ff54007d";
		wait for Clk_period;
		Addr <=  "00000000010100";
		Trees_din <= x"00c1007d";
		wait for Clk_period;
		Addr <=  "00000000010101";
		Trees_din <= x"038a007d";
		wait for Clk_period;
		Addr <=  "00000000010110";
		Trees_din <= x"0615fc0c";
		wait for Clk_period;
		Addr <=  "00000000010111";
		Trees_din <= x"02190304";
		wait for Clk_period;
		Addr <=  "00000000011000";
		Trees_din <= x"03f4007d";
		wait for Clk_period;
		Addr <=  "00000000011001";
		Trees_din <= x"00c00004";
		wait for Clk_period;
		Addr <=  "00000000011010";
		Trees_din <= x"00e2007d";
		wait for Clk_period;
		Addr <=  "00000000011011";
		Trees_din <= x"ff71007d";
		wait for Clk_period;
		Addr <=  "00000000011100";
		Trees_din <= x"0123d704";
		wait for Clk_period;
		Addr <=  "00000000011101";
		Trees_din <= x"ff5e007d";
		wait for Clk_period;
		Addr <=  "00000000011110";
		Trees_din <= x"0203007d";
		wait for Clk_period;
		Addr <=  "00000000011111";
		Trees_din <= x"010e902c";
		wait for Clk_period;
		Addr <=  "00000000100000";
		Trees_din <= x"0105d60c";
		wait for Clk_period;
		Addr <=  "00000000100001";
		Trees_din <= x"0b076904";
		wait for Clk_period;
		Addr <=  "00000000100010";
		Trees_din <= x"ff550111";
		wait for Clk_period;
		Addr <=  "00000000100011";
		Trees_din <= x"12008404";
		wait for Clk_period;
		Addr <=  "00000000100100";
		Trees_din <= x"00340111";
		wait for Clk_period;
		Addr <=  "00000000100101";
		Trees_din <= x"ff710111";
		wait for Clk_period;
		Addr <=  "00000000100110";
		Trees_din <= x"00f56610";
		wait for Clk_period;
		Addr <=  "00000000100111";
		Trees_din <= x"00e76404";
		wait for Clk_period;
		Addr <=  "00000000101000";
		Trees_din <= x"ff570111";
		wait for Clk_period;
		Addr <=  "00000000101001";
		Trees_din <= x"05ffcd04";
		wait for Clk_period;
		Addr <=  "00000000101010";
		Trees_din <= x"ff630111";
		wait for Clk_period;
		Addr <=  "00000000101011";
		Trees_din <= x"0509dd04";
		wait for Clk_period;
		Addr <=  "00000000101100";
		Trees_din <= x"01500111";
		wait for Clk_period;
		Addr <=  "00000000101101";
		Trees_din <= x"ff770111";
		wait for Clk_period;
		Addr <=  "00000000101110";
		Trees_din <= x"020a690c";
		wait for Clk_period;
		Addr <=  "00000000101111";
		Trees_din <= x"06047108";
		wait for Clk_period;
		Addr <=  "00000000110000";
		Trees_din <= x"05075404";
		wait for Clk_period;
		Addr <=  "00000000110001";
		Trees_din <= x"01cc0111";
		wait for Clk_period;
		Addr <=  "00000000110010";
		Trees_din <= x"ffa30111";
		wait for Clk_period;
		Addr <=  "00000000110011";
		Trees_din <= x"ff9d0111";
		wait for Clk_period;
		Addr <=  "00000000110100";
		Trees_din <= x"ff790111";
		wait for Clk_period;
		Addr <=  "00000000110101";
		Trees_din <= x"0615fc18";
		wait for Clk_period;
		Addr <=  "00000000110110";
		Trees_din <= x"02190310";
		wait for Clk_period;
		Addr <=  "00000000110111";
		Trees_din <= x"05150f0c";
		wait for Clk_period;
		Addr <=  "00000000111000";
		Trees_din <= x"01124608";
		wait for Clk_period;
		Addr <=  "00000000111001";
		Trees_din <= x"00e23f04";
		wait for Clk_period;
		Addr <=  "00000000111010";
		Trees_din <= x"ff6e0111";
		wait for Clk_period;
		Addr <=  "00000000111011";
		Trees_din <= x"019c0111";
		wait for Clk_period;
		Addr <=  "00000000111100";
		Trees_din <= x"01af0111";
		wait for Clk_period;
		Addr <=  "00000000111101";
		Trees_din <= x"ff810111";
		wait for Clk_period;
		Addr <=  "00000000111110";
		Trees_din <= x"00c00004";
		wait for Clk_period;
		Addr <=  "00000000111111";
		Trees_din <= x"00b30111";
		wait for Clk_period;
		Addr <=  "00000001000000";
		Trees_din <= x"ff640111";
		wait for Clk_period;
		Addr <=  "00000001000001";
		Trees_din <= x"0123d704";
		wait for Clk_period;
		Addr <=  "00000001000010";
		Trees_din <= x"ff5c0111";
		wait for Clk_period;
		Addr <=  "00000001000011";
		Trees_din <= x"01550111";
		wait for Clk_period;
		Addr <=  "00000001000100";
		Trees_din <= x"010e902c";
		wait for Clk_period;
		Addr <=  "00000001000101";
		Trees_din <= x"0105d60c";
		wait for Clk_period;
		Addr <=  "00000001000110";
		Trees_din <= x"0b076904";
		wait for Clk_period;
		Addr <=  "00000001000111";
		Trees_din <= x"ff5901a5";
		wait for Clk_period;
		Addr <=  "00000001001000";
		Trees_din <= x"1a004804";
		wait for Clk_period;
		Addr <=  "00000001001001";
		Trees_din <= x"ff7901a5";
		wait for Clk_period;
		Addr <=  "00000001001010";
		Trees_din <= x"003d01a5";
		wait for Clk_period;
		Addr <=  "00000001001011";
		Trees_din <= x"00f56610";
		wait for Clk_period;
		Addr <=  "00000001001100";
		Trees_din <= x"00e76404";
		wait for Clk_period;
		Addr <=  "00000001001101";
		Trees_din <= x"ff5c01a5";
		wait for Clk_period;
		Addr <=  "00000001001110";
		Trees_din <= x"010d0408";
		wait for Clk_period;
		Addr <=  "00000001001111";
		Trees_din <= x"0d002d04";
		wait for Clk_period;
		Addr <=  "00000001010000";
		Trees_din <= x"00a401a5";
		wait for Clk_period;
		Addr <=  "00000001010001";
		Trees_din <= x"ff6401a5";
		wait for Clk_period;
		Addr <=  "00000001010010";
		Trees_din <= x"015f01a5";
		wait for Clk_period;
		Addr <=  "00000001010011";
		Trees_din <= x"020a690c";
		wait for Clk_period;
		Addr <=  "00000001010100";
		Trees_din <= x"04040108";
		wait for Clk_period;
		Addr <=  "00000001010101";
		Trees_din <= x"18003104";
		wait for Clk_period;
		Addr <=  "00000001010110";
		Trees_din <= x"ffe701a5";
		wait for Clk_period;
		Addr <=  "00000001010111";
		Trees_din <= x"013d01a5";
		wait for Clk_period;
		Addr <=  "00000001011000";
		Trees_din <= x"ff9f01a5";
		wait for Clk_period;
		Addr <=  "00000001011001";
		Trees_din <= x"ff8201a5";
		wait for Clk_period;
		Addr <=  "00000001011010";
		Trees_din <= x"061cb51c";
		wait for Clk_period;
		Addr <=  "00000001011011";
		Trees_din <= x"021b0614";
		wait for Clk_period;
		Addr <=  "00000001011100";
		Trees_din <= x"05150f10";
		wait for Clk_period;
		Addr <=  "00000001011101";
		Trees_din <= x"01124608";
		wait for Clk_period;
		Addr <=  "00000001011110";
		Trees_din <= x"00e23f04";
		wait for Clk_period;
		Addr <=  "00000001011111";
		Trees_din <= x"ff7001a5";
		wait for Clk_period;
		Addr <=  "00000001100000";
		Trees_din <= x"012501a5";
		wait for Clk_period;
		Addr <=  "00000001100001";
		Trees_din <= x"05f5db04";
		wait for Clk_period;
		Addr <=  "00000001100010";
		Trees_din <= x"001101a5";
		wait for Clk_period;
		Addr <=  "00000001100011";
		Trees_din <= x"013501a5";
		wait for Clk_period;
		Addr <=  "00000001100100";
		Trees_din <= x"ff8301a5";
		wait for Clk_period;
		Addr <=  "00000001100101";
		Trees_din <= x"0ef8d304";
		wait for Clk_period;
		Addr <=  "00000001100110";
		Trees_din <= x"008301a5";
		wait for Clk_period;
		Addr <=  "00000001100111";
		Trees_din <= x"ff6801a5";
		wait for Clk_period;
		Addr <=  "00000001101000";
		Trees_din <= x"ff6301a5";
		wait for Clk_period;
		Addr <=  "00000001101001";
		Trees_din <= x"010db630";
		wait for Clk_period;
		Addr <=  "00000001101010";
		Trees_din <= x"0105d60c";
		wait for Clk_period;
		Addr <=  "00000001101011";
		Trees_din <= x"0b076904";
		wait for Clk_period;
		Addr <=  "00000001101100";
		Trees_din <= x"ff5d0249";
		wait for Clk_period;
		Addr <=  "00000001101101";
		Trees_din <= x"09fcb804";
		wait for Clk_period;
		Addr <=  "00000001101110";
		Trees_din <= x"00450249";
		wait for Clk_period;
		Addr <=  "00000001101111";
		Trees_din <= x"ff800249";
		wait for Clk_period;
		Addr <=  "00000001110000";
		Trees_din <= x"00f56610";
		wait for Clk_period;
		Addr <=  "00000001110001";
		Trees_din <= x"0d002d08";
		wait for Clk_period;
		Addr <=  "00000001110010";
		Trees_din <= x"1a004504";
		wait for Clk_period;
		Addr <=  "00000001110011";
		Trees_din <= x"00bf0249";
		wait for Clk_period;
		Addr <=  "00000001110100";
		Trees_din <= x"ff910249";
		wait for Clk_period;
		Addr <=  "00000001110101";
		Trees_din <= x"1b03d704";
		wait for Clk_period;
		Addr <=  "00000001110110";
		Trees_din <= x"ff5f0249";
		wait for Clk_period;
		Addr <=  "00000001110111";
		Trees_din <= x"00010249";
		wait for Clk_period;
		Addr <=  "00000001111000";
		Trees_din <= x"020a6910";
		wait for Clk_period;
		Addr <=  "00000001111001";
		Trees_din <= x"02ff3808";
		wait for Clk_period;
		Addr <=  "00000001111010";
		Trees_din <= x"0d00b604";
		wait for Clk_period;
		Addr <=  "00000001111011";
		Trees_din <= x"00140249";
		wait for Clk_period;
		Addr <=  "00000001111100";
		Trees_din <= x"ff9b0249";
		wait for Clk_period;
		Addr <=  "00000001111101";
		Trees_din <= x"18003104";
		wait for Clk_period;
		Addr <=  "00000001111110";
		Trees_din <= x"fffa0249";
		wait for Clk_period;
		Addr <=  "00000001111111";
		Trees_din <= x"00f80249";
		wait for Clk_period;
		Addr <=  "00000010000000";
		Trees_din <= x"ff8c0249";
		wait for Clk_period;
		Addr <=  "00000010000001";
		Trees_din <= x"0615fc1c";
		wait for Clk_period;
		Addr <=  "00000010000010";
		Trees_din <= x"02186814";
		wait for Clk_period;
		Addr <=  "00000010000011";
		Trees_din <= x"05150f10";
		wait for Clk_period;
		Addr <=  "00000010000100";
		Trees_din <= x"05f5db08";
		wait for Clk_period;
		Addr <=  "00000010000101";
		Trees_din <= x"18003904";
		wait for Clk_period;
		Addr <=  "00000010000110";
		Trees_din <= x"ff7b0249";
		wait for Clk_period;
		Addr <=  "00000010000111";
		Trees_din <= x"00ae0249";
		wait for Clk_period;
		Addr <=  "00000010001000";
		Trees_din <= x"04171604";
		wait for Clk_period;
		Addr <=  "00000010001001";
		Trees_din <= x"00f90249";
		wait for Clk_period;
		Addr <=  "00000010001010";
		Trees_din <= x"00770249";
		wait for Clk_period;
		Addr <=  "00000010001011";
		Trees_din <= x"ff930249";
		wait for Clk_period;
		Addr <=  "00000010001100";
		Trees_din <= x"012a7d04";
		wait for Clk_period;
		Addr <=  "00000010001101";
		Trees_din <= x"ff680249";
		wait for Clk_period;
		Addr <=  "00000010001110";
		Trees_din <= x"010f0249";
		wait for Clk_period;
		Addr <=  "00000010001111";
		Trees_din <= x"0123d704";
		wait for Clk_period;
		Addr <=  "00000010010000";
		Trees_din <= x"ff660249";
		wait for Clk_period;
		Addr <=  "00000010010001";
		Trees_din <= x"00c80249";
		wait for Clk_period;
		Addr <=  "00000010010010";
		Trees_din <= x"010db630";
		wait for Clk_period;
		Addr <=  "00000010010011";
		Trees_din <= x"0105190c";
		wait for Clk_period;
		Addr <=  "00000010010100";
		Trees_din <= x"0b076904";
		wait for Clk_period;
		Addr <=  "00000010010101";
		Trees_din <= x"ff5f02d5";
		wait for Clk_period;
		Addr <=  "00000010010110";
		Trees_din <= x"11003904";
		wait for Clk_period;
		Addr <=  "00000010010111";
		Trees_din <= x"004702d5";
		wait for Clk_period;
		Addr <=  "00000010011000";
		Trees_din <= x"ff8902d5";
		wait for Clk_period;
		Addr <=  "00000010011001";
		Trees_din <= x"00f56610";
		wait for Clk_period;
		Addr <=  "00000010011010";
		Trees_din <= x"0d002d08";
		wait for Clk_period;
		Addr <=  "00000010011011";
		Trees_din <= x"18003704";
		wait for Clk_period;
		Addr <=  "00000010011100";
		Trees_din <= x"00b302d5";
		wait for Clk_period;
		Addr <=  "00000010011101";
		Trees_din <= x"ff9302d5";
		wait for Clk_period;
		Addr <=  "00000010011110";
		Trees_din <= x"0f04b704";
		wait for Clk_period;
		Addr <=  "00000010011111";
		Trees_din <= x"ff6202d5";
		wait for Clk_period;
		Addr <=  "00000010100000";
		Trees_din <= x"000602d5";
		wait for Clk_period;
		Addr <=  "00000010100001";
		Trees_din <= x"020a6910";
		wait for Clk_period;
		Addr <=  "00000010100010";
		Trees_din <= x"1a003f08";
		wait for Clk_period;
		Addr <=  "00000010100011";
		Trees_din <= x"0b011704";
		wait for Clk_period;
		Addr <=  "00000010100100";
		Trees_din <= x"006602d5";
		wait for Clk_period;
		Addr <=  "00000010100101";
		Trees_din <= x"ff7f02d5";
		wait for Clk_period;
		Addr <=  "00000010100110";
		Trees_din <= x"0bfc2e04";
		wait for Clk_period;
		Addr <=  "00000010100111";
		Trees_din <= x"004102d5";
		wait for Clk_period;
		Addr <=  "00000010101000";
		Trees_din <= x"00ed02d5";
		wait for Clk_period;
		Addr <=  "00000010101001";
		Trees_din <= x"ff8902d5";
		wait for Clk_period;
		Addr <=  "00000010101010";
		Trees_din <= x"061cb514";
		wait for Clk_period;
		Addr <=  "00000010101011";
		Trees_din <= x"021cf410";
		wait for Clk_period;
		Addr <=  "00000010101100";
		Trees_din <= x"0118430c";
		wait for Clk_period;
		Addr <=  "00000010101101";
		Trees_din <= x"060d1808";
		wait for Clk_period;
		Addr <=  "00000010101110";
		Trees_din <= x"00ce5b04";
		wait for Clk_period;
		Addr <=  "00000010101111";
		Trees_din <= x"ffd402d5";
		wait for Clk_period;
		Addr <=  "00000010110000";
		Trees_din <= x"00db02d5";
		wait for Clk_period;
		Addr <=  "00000010110001";
		Trees_din <= x"ff5b02d5";
		wait for Clk_period;
		Addr <=  "00000010110010";
		Trees_din <= x"00e002d5";
		wait for Clk_period;
		Addr <=  "00000010110011";
		Trees_din <= x"ff7202d5";
		wait for Clk_period;
		Addr <=  "00000010110100";
		Trees_din <= x"ff6d02d5";
		wait for Clk_period;
		Addr <=  "00000010110101";
		Trees_din <= x"010db630";
		wait for Clk_period;
		Addr <=  "00000010110110";
		Trees_din <= x"0105190c";
		wait for Clk_period;
		Addr <=  "00000010110111";
		Trees_din <= x"0b076904";
		wait for Clk_period;
		Addr <=  "00000010111000";
		Trees_din <= x"ff620369";
		wait for Clk_period;
		Addr <=  "00000010111001";
		Trees_din <= x"14002504";
		wait for Clk_period;
		Addr <=  "00000010111010";
		Trees_din <= x"00470369";
		wait for Clk_period;
		Addr <=  "00000010111011";
		Trees_din <= x"ff920369";
		wait for Clk_period;
		Addr <=  "00000010111100";
		Trees_din <= x"00f56610";
		wait for Clk_period;
		Addr <=  "00000010111101";
		Trees_din <= x"0d002d08";
		wait for Clk_period;
		Addr <=  "00000010111110";
		Trees_din <= x"00e9ab04";
		wait for Clk_period;
		Addr <=  "00000010111111";
		Trees_din <= x"ff9c0369";
		wait for Clk_period;
		Addr <=  "00000011000000";
		Trees_din <= x"00990369";
		wait for Clk_period;
		Addr <=  "00000011000001";
		Trees_din <= x"1b03d704";
		wait for Clk_period;
		Addr <=  "00000011000010";
		Trees_din <= x"ff650369";
		wait for Clk_period;
		Addr <=  "00000011000011";
		Trees_din <= x"000d0369";
		wait for Clk_period;
		Addr <=  "00000011000100";
		Trees_din <= x"020a6910";
		wait for Clk_period;
		Addr <=  "00000011000101";
		Trees_din <= x"0c014008";
		wait for Clk_period;
		Addr <=  "00000011000110";
		Trees_din <= x"1a003e04";
		wait for Clk_period;
		Addr <=  "00000011000111";
		Trees_din <= x"00290369";
		wait for Clk_period;
		Addr <=  "00000011001000";
		Trees_din <= x"00cc0369";
		wait for Clk_period;
		Addr <=  "00000011001001";
		Trees_din <= x"01096504";
		wait for Clk_period;
		Addr <=  "00000011001010";
		Trees_din <= x"ffa80369";
		wait for Clk_period;
		Addr <=  "00000011001011";
		Trees_din <= x"00720369";
		wait for Clk_period;
		Addr <=  "00000011001100";
		Trees_din <= x"ff920369";
		wait for Clk_period;
		Addr <=  "00000011001101";
		Trees_din <= x"061cb518";
		wait for Clk_period;
		Addr <=  "00000011001110";
		Trees_din <= x"021bef10";
		wait for Clk_period;
		Addr <=  "00000011001111";
		Trees_din <= x"05150f0c";
		wait for Clk_period;
		Addr <=  "00000011010000";
		Trees_din <= x"01184308";
		wait for Clk_period;
		Addr <=  "00000011010001";
		Trees_din <= x"060d1804";
		wait for Clk_period;
		Addr <=  "00000011010010";
		Trees_din <= x"00a80369";
		wait for Clk_period;
		Addr <=  "00000011010011";
		Trees_din <= x"ff670369";
		wait for Clk_period;
		Addr <=  "00000011010100";
		Trees_din <= x"00ca0369";
		wait for Clk_period;
		Addr <=  "00000011010101";
		Trees_din <= x"ff960369";
		wait for Clk_period;
		Addr <=  "00000011010110";
		Trees_din <= x"030b9804";
		wait for Clk_period;
		Addr <=  "00000011010111";
		Trees_din <= x"ff780369";
		wait for Clk_period;
		Addr <=  "00000011011000";
		Trees_din <= x"00260369";
		wait for Clk_period;
		Addr <=  "00000011011001";
		Trees_din <= x"ff730369";
		wait for Clk_period;
		Addr <=  "00000011011010";
		Trees_din <= x"010d0438";
		wait for Clk_period;
		Addr <=  "00000011011011";
		Trees_din <= x"01051914";
		wait for Clk_period;
		Addr <=  "00000011011100";
		Trees_din <= x"0b07690c";
		wait for Clk_period;
		Addr <=  "00000011011101";
		Trees_din <= x"0ffb1c08";
		wait for Clk_period;
		Addr <=  "00000011011110";
		Trees_din <= x"0a00a604";
		wait for Clk_period;
		Addr <=  "00000011011111";
		Trees_din <= x"00470415";
		wait for Clk_period;
		Addr <=  "00000011100000";
		Trees_din <= x"ff7a0415";
		wait for Clk_period;
		Addr <=  "00000011100001";
		Trees_din <= x"ff630415";
		wait for Clk_period;
		Addr <=  "00000011100010";
		Trees_din <= x"03fdbf04";
		wait for Clk_period;
		Addr <=  "00000011100011";
		Trees_din <= x"00480415";
		wait for Clk_period;
		Addr <=  "00000011100100";
		Trees_din <= x"ff9c0415";
		wait for Clk_period;
		Addr <=  "00000011100101";
		Trees_din <= x"00f5660c";
		wait for Clk_period;
		Addr <=  "00000011100110";
		Trees_din <= x"0d002d08";
		wait for Clk_period;
		Addr <=  "00000011100111";
		Trees_din <= x"01096504";
		wait for Clk_period;
		Addr <=  "00000011101000";
		Trees_din <= x"ffa60415";
		wait for Clk_period;
		Addr <=  "00000011101001";
		Trees_din <= x"008c0415";
		wait for Clk_period;
		Addr <=  "00000011101010";
		Trees_din <= x"ff680415";
		wait for Clk_period;
		Addr <=  "00000011101011";
		Trees_din <= x"0c01400c";
		wait for Clk_period;
		Addr <=  "00000011101100";
		Trees_din <= x"1a003e04";
		wait for Clk_period;
		Addr <=  "00000011101101";
		Trees_din <= x"00040415";
		wait for Clk_period;
		Addr <=  "00000011101110";
		Trees_din <= x"14006904";
		wait for Clk_period;
		Addr <=  "00000011101111";
		Trees_din <= x"00390415";
		wait for Clk_period;
		Addr <=  "00000011110000";
		Trees_din <= x"00b10415";
		wait for Clk_period;
		Addr <=  "00000011110001";
		Trees_din <= x"16000008";
		wait for Clk_period;
		Addr <=  "00000011110010";
		Trees_din <= x"08005304";
		wait for Clk_period;
		Addr <=  "00000011110011";
		Trees_din <= x"00600415";
		wait for Clk_period;
		Addr <=  "00000011110100";
		Trees_din <= x"fff20415";
		wait for Clk_period;
		Addr <=  "00000011110101";
		Trees_din <= x"ff7d0415";
		wait for Clk_period;
		Addr <=  "00000011110110";
		Trees_din <= x"061cb51c";
		wait for Clk_period;
		Addr <=  "00000011110111";
		Trees_din <= x"0217b314";
		wait for Clk_period;
		Addr <=  "00000011111000";
		Trees_din <= x"0614d40c";
		wait for Clk_period;
		Addr <=  "00000011111001";
		Trees_din <= x"0513e608";
		wait for Clk_period;
		Addr <=  "00000011111010";
		Trees_din <= x"04121004";
		wait for Clk_period;
		Addr <=  "00000011111011";
		Trees_din <= x"00b70415";
		wait for Clk_period;
		Addr <=  "00000011111100";
		Trees_din <= x"00430415";
		wait for Clk_period;
		Addr <=  "00000011111101";
		Trees_din <= x"ffa50415";
		wait for Clk_period;
		Addr <=  "00000011111110";
		Trees_din <= x"011fa004";
		wait for Clk_period;
		Addr <=  "00000011111111";
		Trees_din <= x"ff800415";
		wait for Clk_period;
		Addr <=  "00000100000000";
		Trees_din <= x"009e0415";
		wait for Clk_period;
		Addr <=  "00000100000001";
		Trees_din <= x"012a7d04";
		wait for Clk_period;
		Addr <=  "00000100000010";
		Trees_din <= x"ff700415";
		wait for Clk_period;
		Addr <=  "00000100000011";
		Trees_din <= x"00af0415";
		wait for Clk_period;
		Addr <=  "00000100000100";
		Trees_din <= x"ff780415";
		wait for Clk_period;
		Addr <=  "00000100000101";
		Trees_din <= x"01096524";
		wait for Clk_period;
		Addr <=  "00000100000110";
		Trees_din <= x"0105190c";
		wait for Clk_period;
		Addr <=  "00000100000111";
		Trees_din <= x"10fc6f08";
		wait for Clk_period;
		Addr <=  "00000100001000";
		Trees_din <= x"19008204";
		wait for Clk_period;
		Addr <=  "00000100001001";
		Trees_din <= x"00e004a1";
		wait for Clk_period;
		Addr <=  "00000100001010";
		Trees_din <= x"ff7704a1";
		wait for Clk_period;
		Addr <=  "00000100001011";
		Trees_din <= x"ff6404a1";
		wait for Clk_period;
		Addr <=  "00000100001100";
		Trees_din <= x"00fdf110";
		wait for Clk_period;
		Addr <=  "00000100001101";
		Trees_din <= x"00f95f08";
		wait for Clk_period;
		Addr <=  "00000100001110";
		Trees_din <= x"12007d04";
		wait for Clk_period;
		Addr <=  "00000100001111";
		Trees_din <= x"fffa04a1";
		wait for Clk_period;
		Addr <=  "00000100010000";
		Trees_din <= x"ff6d04a1";
		wait for Clk_period;
		Addr <=  "00000100010001";
		Trees_din <= x"17004104";
		wait for Clk_period;
		Addr <=  "00000100010010";
		Trees_din <= x"ff9104a1";
		wait for Clk_period;
		Addr <=  "00000100010011";
		Trees_din <= x"003c04a1";
		wait for Clk_period;
		Addr <=  "00000100010100";
		Trees_din <= x"06fe6f04";
		wait for Clk_period;
		Addr <=  "00000100010101";
		Trees_din <= x"001204a1";
		wait for Clk_period;
		Addr <=  "00000100010110";
		Trees_din <= x"00a404a1";
		wait for Clk_period;
		Addr <=  "00000100010111";
		Trees_din <= x"0615fc1c";
		wait for Clk_period;
		Addr <=  "00000100011000";
		Trees_din <= x"0216d914";
		wait for Clk_period;
		Addr <=  "00000100011001";
		Trees_din <= x"0513e610";
		wait for Clk_period;
		Addr <=  "00000100011010";
		Trees_din <= x"01124608";
		wait for Clk_period;
		Addr <=  "00000100011011";
		Trees_din <= x"00e23f04";
		wait for Clk_period;
		Addr <=  "00000100011100";
		Trees_din <= x"ff7a04a1";
		wait for Clk_period;
		Addr <=  "00000100011101";
		Trees_din <= x"009604a1";
		wait for Clk_period;
		Addr <=  "00000100011110";
		Trees_din <= x"05f5db04";
		wait for Clk_period;
		Addr <=  "00000100011111";
		Trees_din <= x"fffa04a1";
		wait for Clk_period;
		Addr <=  "00000100100000";
		Trees_din <= x"00a904a1";
		wait for Clk_period;
		Addr <=  "00000100100001";
		Trees_din <= x"ffb104a1";
		wait for Clk_period;
		Addr <=  "00000100100010";
		Trees_din <= x"012a7d04";
		wait for Clk_period;
		Addr <=  "00000100100011";
		Trees_din <= x"ff7304a1";
		wait for Clk_period;
		Addr <=  "00000100100100";
		Trees_din <= x"009804a1";
		wait for Clk_period;
		Addr <=  "00000100100101";
		Trees_din <= x"0123d704";
		wait for Clk_period;
		Addr <=  "00000100100110";
		Trees_din <= x"ff7404a1";
		wait for Clk_period;
		Addr <=  "00000100100111";
		Trees_din <= x"006b04a1";
		wait for Clk_period;
		Addr <=  "00000100101000";
		Trees_din <= x"0109652c";
		wait for Clk_period;
		Addr <=  "00000100101001";
		Trees_din <= x"01051914";
		wait for Clk_period;
		Addr <=  "00000100101010";
		Trees_din <= x"10fc6f08";
		wait for Clk_period;
		Addr <=  "00000100101011";
		Trees_din <= x"1a004f04";
		wait for Clk_period;
		Addr <=  "00000100101100";
		Trees_din <= x"ff7c0545";
		wait for Clk_period;
		Addr <=  "00000100101101";
		Trees_din <= x"00da0545";
		wait for Clk_period;
		Addr <=  "00000100101110";
		Trees_din <= x"0ef83c08";
		wait for Clk_period;
		Addr <=  "00000100101111";
		Trees_din <= x"0506ce04";
		wait for Clk_period;
		Addr <=  "00000100110000";
		Trees_din <= x"ff7d0545";
		wait for Clk_period;
		Addr <=  "00000100110001";
		Trees_din <= x"00400545";
		wait for Clk_period;
		Addr <=  "00000100110010";
		Trees_din <= x"ff640545";
		wait for Clk_period;
		Addr <=  "00000100110011";
		Trees_din <= x"00fdf110";
		wait for Clk_period;
		Addr <=  "00000100110100";
		Trees_din <= x"06fe4108";
		wait for Clk_period;
		Addr <=  "00000100110101";
		Trees_din <= x"10022904";
		wait for Clk_period;
		Addr <=  "00000100110110";
		Trees_din <= x"ffa50545";
		wait for Clk_period;
		Addr <=  "00000100110111";
		Trees_din <= x"00180545";
		wait for Clk_period;
		Addr <=  "00000100111000";
		Trees_din <= x"02fb8e04";
		wait for Clk_period;
		Addr <=  "00000100111001";
		Trees_din <= x"ffea0545";
		wait for Clk_period;
		Addr <=  "00000100111010";
		Trees_din <= x"ff6e0545";
		wait for Clk_period;
		Addr <=  "00000100111011";
		Trees_din <= x"1b011604";
		wait for Clk_period;
		Addr <=  "00000100111100";
		Trees_din <= x"008b0545";
		wait for Clk_period;
		Addr <=  "00000100111101";
		Trees_din <= x"00200545";
		wait for Clk_period;
		Addr <=  "00000100111110";
		Trees_din <= x"01184320";
		wait for Clk_period;
		Addr <=  "00000100111111";
		Trees_din <= x"00d71810";
		wait for Clk_period;
		Addr <=  "00000101000000";
		Trees_din <= x"01152c04";
		wait for Clk_period;
		Addr <=  "00000101000001";
		Trees_din <= x"ff6d0545";
		wait for Clk_period;
		Addr <=  "00000101000010";
		Trees_din <= x"060c5d08";
		wait for Clk_period;
		Addr <=  "00000101000011";
		Trees_din <= x"15024d04";
		wait for Clk_period;
		Addr <=  "00000101000100";
		Trees_din <= x"00690545";
		wait for Clk_period;
		Addr <=  "00000101000101";
		Trees_din <= x"000c0545";
		wait for Clk_period;
		Addr <=  "00000101000110";
		Trees_din <= x"ff8b0545";
		wait for Clk_period;
		Addr <=  "00000101000111";
		Trees_din <= x"060af00c";
		wait for Clk_period;
		Addr <=  "00000101001000";
		Trees_din <= x"05085508";
		wait for Clk_period;
		Addr <=  "00000101001001";
		Trees_din <= x"05f5db04";
		wait for Clk_period;
		Addr <=  "00000101001010";
		Trees_din <= x"fffe0545";
		wait for Clk_period;
		Addr <=  "00000101001011";
		Trees_din <= x"009e0545";
		wait for Clk_period;
		Addr <=  "00000101001100";
		Trees_din <= x"fffb0545";
		wait for Clk_period;
		Addr <=  "00000101001101";
		Trees_din <= x"ffa20545";
		wait for Clk_period;
		Addr <=  "00000101001110";
		Trees_din <= x"061cb504";
		wait for Clk_period;
		Addr <=  "00000101001111";
		Trees_din <= x"009f0545";
		wait for Clk_period;
		Addr <=  "00000101010000";
		Trees_din <= x"ffa70545";
		wait for Clk_period;
		Addr <=  "00000101010001";
		Trees_din <= x"0109652c";
		wait for Clk_period;
		Addr <=  "00000101010010";
		Trees_din <= x"01051914";
		wait for Clk_period;
		Addr <=  "00000101010011";
		Trees_din <= x"10fc6f08";
		wait for Clk_period;
		Addr <=  "00000101010100";
		Trees_din <= x"1a005104";
		wait for Clk_period;
		Addr <=  "00000101010101";
		Trees_din <= x"ff8205f9";
		wait for Clk_period;
		Addr <=  "00000101010110";
		Trees_din <= x"00ca05f9";
		wait for Clk_period;
		Addr <=  "00000101010111";
		Trees_din <= x"0ef83c08";
		wait for Clk_period;
		Addr <=  "00000101011000";
		Trees_din <= x"07005404";
		wait for Clk_period;
		Addr <=  "00000101011001";
		Trees_din <= x"004a05f9";
		wait for Clk_period;
		Addr <=  "00000101011010";
		Trees_din <= x"ff8305f9";
		wait for Clk_period;
		Addr <=  "00000101011011";
		Trees_din <= x"ff6505f9";
		wait for Clk_period;
		Addr <=  "00000101011100";
		Trees_din <= x"00fdf110";
		wait for Clk_period;
		Addr <=  "00000101011101";
		Trees_din <= x"06fe4108";
		wait for Clk_period;
		Addr <=  "00000101011110";
		Trees_din <= x"06fc9b04";
		wait for Clk_period;
		Addr <=  "00000101011111";
		Trees_din <= x"ffad05f9";
		wait for Clk_period;
		Addr <=  "00000101100000";
		Trees_din <= x"001705f9";
		wait for Clk_period;
		Addr <=  "00000101100001";
		Trees_din <= x"1c002604";
		wait for Clk_period;
		Addr <=  "00000101100010";
		Trees_din <= x"ffe805f9";
		wait for Clk_period;
		Addr <=  "00000101100011";
		Trees_din <= x"ff7205f9";
		wait for Clk_period;
		Addr <=  "00000101100100";
		Trees_din <= x"03fcaf04";
		wait for Clk_period;
		Addr <=  "00000101100101";
		Trees_din <= x"002405f9";
		wait for Clk_period;
		Addr <=  "00000101100110";
		Trees_din <= x"007f05f9";
		wait for Clk_period;
		Addr <=  "00000101100111";
		Trees_din <= x"01184320";
		wait for Clk_period;
		Addr <=  "00000101101000";
		Trees_din <= x"00d71810";
		wait for Clk_period;
		Addr <=  "00000101101001";
		Trees_din <= x"01152c04";
		wait for Clk_period;
		Addr <=  "00000101101010";
		Trees_din <= x"ff7105f9";
		wait for Clk_period;
		Addr <=  "00000101101011";
		Trees_din <= x"060c5d08";
		wait for Clk_period;
		Addr <=  "00000101101100";
		Trees_din <= x"020bd204";
		wait for Clk_period;
		Addr <=  "00000101101101";
		Trees_din <= x"005e05f9";
		wait for Clk_period;
		Addr <=  "00000101101110";
		Trees_din <= x"001105f9";
		wait for Clk_period;
		Addr <=  "00000101101111";
		Trees_din <= x"ff9505f9";
		wait for Clk_period;
		Addr <=  "00000101110000";
		Trees_din <= x"060af00c";
		wait for Clk_period;
		Addr <=  "00000101110001";
		Trees_din <= x"00e5d908";
		wait for Clk_period;
		Addr <=  "00000101110010";
		Trees_din <= x"010f7504";
		wait for Clk_period;
		Addr <=  "00000101110011";
		Trees_din <= x"ff9e05f9";
		wait for Clk_period;
		Addr <=  "00000101110100";
		Trees_din <= x"007d05f9";
		wait for Clk_period;
		Addr <=  "00000101110101";
		Trees_din <= x"009905f9";
		wait for Clk_period;
		Addr <=  "00000101110110";
		Trees_din <= x"ffae05f9";
		wait for Clk_period;
		Addr <=  "00000101110111";
		Trees_din <= x"061cb50c";
		wait for Clk_period;
		Addr <=  "00000101111000";
		Trees_din <= x"07004d04";
		wait for Clk_period;
		Addr <=  "00000101111001";
		Trees_din <= x"002c05f9";
		wait for Clk_period;
		Addr <=  "00000101111010";
		Trees_din <= x"0615fc04";
		wait for Clk_period;
		Addr <=  "00000101111011";
		Trees_din <= x"009d05f9";
		wait for Clk_period;
		Addr <=  "00000101111100";
		Trees_din <= x"004005f9";
		wait for Clk_period;
		Addr <=  "00000101111101";
		Trees_din <= x"ffad05f9";
		wait for Clk_period;
		Addr <=  "00000101111110";
		Trees_din <= x"01096528";
		wait for Clk_period;
		Addr <=  "00000101111111";
		Trees_din <= x"01051914";
		wait for Clk_period;
		Addr <=  "00000110000000";
		Trees_din <= x"10fc6f08";
		wait for Clk_period;
		Addr <=  "00000110000001";
		Trees_din <= x"1a005104";
		wait for Clk_period;
		Addr <=  "00000110000010";
		Trees_din <= x"ff89067d";
		wait for Clk_period;
		Addr <=  "00000110000011";
		Trees_din <= x"00aa067d";
		wait for Clk_period;
		Addr <=  "00000110000100";
		Trees_din <= x"0ef83c08";
		wait for Clk_period;
		Addr <=  "00000110000101";
		Trees_din <= x"04fe8b04";
		wait for Clk_period;
		Addr <=  "00000110000110";
		Trees_din <= x"0040067d";
		wait for Clk_period;
		Addr <=  "00000110000111";
		Trees_din <= x"ff8b067d";
		wait for Clk_period;
		Addr <=  "00000110001000";
		Trees_din <= x"ff66067d";
		wait for Clk_period;
		Addr <=  "00000110001001";
		Trees_din <= x"00fdf110";
		wait for Clk_period;
		Addr <=  "00000110001010";
		Trees_din <= x"06fe4108";
		wait for Clk_period;
		Addr <=  "00000110001011";
		Trees_din <= x"03fbeb04";
		wait for Clk_period;
		Addr <=  "00000110001100";
		Trees_din <= x"ffc2067d";
		wait for Clk_period;
		Addr <=  "00000110001101";
		Trees_din <= x"0017067d";
		wait for Clk_period;
		Addr <=  "00000110001110";
		Trees_din <= x"07005b04";
		wait for Clk_period;
		Addr <=  "00000110001111";
		Trees_din <= x"ff77067d";
		wait for Clk_period;
		Addr <=  "00000110010000";
		Trees_din <= x"ffe5067d";
		wait for Clk_period;
		Addr <=  "00000110010001";
		Trees_din <= x"0060067d";
		wait for Clk_period;
		Addr <=  "00000110010010";
		Trees_din <= x"021a0314";
		wait for Clk_period;
		Addr <=  "00000110010011";
		Trees_din <= x"061cb510";
		wait for Clk_period;
		Addr <=  "00000110010100";
		Trees_din <= x"0118430c";
		wait for Clk_period;
		Addr <=  "00000110010101";
		Trees_din <= x"060d1808";
		wait for Clk_period;
		Addr <=  "00000110010110";
		Trees_din <= x"04078904";
		wait for Clk_period;
		Addr <=  "00000110010111";
		Trees_din <= x"007e067d";
		wait for Clk_period;
		Addr <=  "00000110011000";
		Trees_din <= x"ffed067d";
		wait for Clk_period;
		Addr <=  "00000110011001";
		Trees_din <= x"ff83067d";
		wait for Clk_period;
		Addr <=  "00000110011010";
		Trees_din <= x"009b067d";
		wait for Clk_period;
		Addr <=  "00000110011011";
		Trees_din <= x"ff8f067d";
		wait for Clk_period;
		Addr <=  "00000110011100";
		Trees_din <= x"1403ae04";
		wait for Clk_period;
		Addr <=  "00000110011101";
		Trees_din <= x"ff85067d";
		wait for Clk_period;
		Addr <=  "00000110011110";
		Trees_din <= x"0016067d";
		wait for Clk_period;
		Addr <=  "00000110011111";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00000110100000";
		Trees_din <= x"01081b20";
		wait for Clk_period;
		Addr <=  "00000110100001";
		Trees_din <= x"10fc6f08";
		wait for Clk_period;
		Addr <=  "00000110100010";
		Trees_din <= x"1a005104";
		wait for Clk_period;
		Addr <=  "00000110100011";
		Trees_din <= x"ff910725";
		wait for Clk_period;
		Addr <=  "00000110100100";
		Trees_din <= x"00910725";
		wait for Clk_period;
		Addr <=  "00000110100101";
		Trees_din <= x"0105190c";
		wait for Clk_period;
		Addr <=  "00000110100110";
		Trees_din <= x"0ef83c08";
		wait for Clk_period;
		Addr <=  "00000110100111";
		Trees_din <= x"0d019704";
		wait for Clk_period;
		Addr <=  "00000110101000";
		Trees_din <= x"ff920725";
		wait for Clk_period;
		Addr <=  "00000110101001";
		Trees_din <= x"00490725";
		wait for Clk_period;
		Addr <=  "00000110101010";
		Trees_din <= x"ff670725";
		wait for Clk_period;
		Addr <=  "00000110101011";
		Trees_din <= x"00fdf108";
		wait for Clk_period;
		Addr <=  "00000110101100";
		Trees_din <= x"06fd1a04";
		wait for Clk_period;
		Addr <=  "00000110101101";
		Trees_din <= x"ffed0725";
		wait for Clk_period;
		Addr <=  "00000110101110";
		Trees_din <= x"ff820725";
		wait for Clk_period;
		Addr <=  "00000110101111";
		Trees_din <= x"00530725";
		wait for Clk_period;
		Addr <=  "00000110110000";
		Trees_din <= x"0116f124";
		wait for Clk_period;
		Addr <=  "00000110110001";
		Trees_din <= x"00e5d914";
		wait for Clk_period;
		Addr <=  "00000110110010";
		Trees_din <= x"01124608";
		wait for Clk_period;
		Addr <=  "00000110110011";
		Trees_din <= x"0601fd04";
		wait for Clk_period;
		Addr <=  "00000110110100";
		Trees_din <= x"ffda0725";
		wait for Clk_period;
		Addr <=  "00000110110101";
		Trees_din <= x"ff790725";
		wait for Clk_period;
		Addr <=  "00000110110110";
		Trees_din <= x"00d25d04";
		wait for Clk_period;
		Addr <=  "00000110110111";
		Trees_din <= x"ffa10725";
		wait for Clk_period;
		Addr <=  "00000110111000";
		Trees_din <= x"0a013704";
		wait for Clk_period;
		Addr <=  "00000110111001";
		Trees_din <= x"006c0725";
		wait for Clk_period;
		Addr <=  "00000110111010";
		Trees_din <= x"00150725";
		wait for Clk_period;
		Addr <=  "00000110111011";
		Trees_din <= x"010d040c";
		wait for Clk_period;
		Addr <=  "00000110111100";
		Trees_din <= x"0efdf604";
		wait for Clk_period;
		Addr <=  "00000110111101";
		Trees_din <= x"006d0725";
		wait for Clk_period;
		Addr <=  "00000110111110";
		Trees_din <= x"0f026a04";
		wait for Clk_period;
		Addr <=  "00000110111111";
		Trees_din <= x"ffa00725";
		wait for Clk_period;
		Addr <=  "00000111000000";
		Trees_din <= x"000b0725";
		wait for Clk_period;
		Addr <=  "00000111000001";
		Trees_din <= x"00910725";
		wait for Clk_period;
		Addr <=  "00000111000010";
		Trees_din <= x"050fb30c";
		wait for Clk_period;
		Addr <=  "00000111000011";
		Trees_din <= x"01184308";
		wait for Clk_period;
		Addr <=  "00000111000100";
		Trees_din <= x"03010304";
		wait for Clk_period;
		Addr <=  "00000111000101";
		Trees_din <= x"00660725";
		wait for Clk_period;
		Addr <=  "00000111000110";
		Trees_din <= x"fff70725";
		wait for Clk_period;
		Addr <=  "00000111000111";
		Trees_din <= x"00880725";
		wait for Clk_period;
		Addr <=  "00000111001000";
		Trees_din <= x"ffd90725";
		wait for Clk_period;
		Addr <=  "00000111001001";
		Trees_din <= x"01081b1c";
		wait for Clk_period;
		Addr <=  "00000111001010";
		Trees_din <= x"10fc6f08";
		wait for Clk_period;
		Addr <=  "00000111001011";
		Trees_din <= x"1a005104";
		wait for Clk_period;
		Addr <=  "00000111001100";
		Trees_din <= x"ff9907a9";
		wait for Clk_period;
		Addr <=  "00000111001101";
		Trees_din <= x"007d07a9";
		wait for Clk_period;
		Addr <=  "00000111001110";
		Trees_din <= x"0105190c";
		wait for Clk_period;
		Addr <=  "00000111001111";
		Trees_din <= x"0ef83c08";
		wait for Clk_period;
		Addr <=  "00000111010000";
		Trees_din <= x"0c038604";
		wait for Clk_period;
		Addr <=  "00000111010001";
		Trees_din <= x"ff9a07a9";
		wait for Clk_period;
		Addr <=  "00000111010010";
		Trees_din <= x"004607a9";
		wait for Clk_period;
		Addr <=  "00000111010011";
		Trees_din <= x"ff6707a9";
		wait for Clk_period;
		Addr <=  "00000111010100";
		Trees_din <= x"00f95f04";
		wait for Clk_period;
		Addr <=  "00000111010101";
		Trees_din <= x"ff8807a9";
		wait for Clk_period;
		Addr <=  "00000111010110";
		Trees_din <= x"002e07a9";
		wait for Clk_period;
		Addr <=  "00000111010111";
		Trees_din <= x"021a0320";
		wait for Clk_period;
		Addr <=  "00000111011000";
		Trees_din <= x"061cb51c";
		wait for Clk_period;
		Addr <=  "00000111011001";
		Trees_din <= x"0112460c";
		wait for Clk_period;
		Addr <=  "00000111011010";
		Trees_din <= x"00e5d904";
		wait for Clk_period;
		Addr <=  "00000111011011";
		Trees_din <= x"ff9807a9";
		wait for Clk_period;
		Addr <=  "00000111011100";
		Trees_din <= x"15f9bc04";
		wait for Clk_period;
		Addr <=  "00000111011101";
		Trees_din <= x"ffea07a9";
		wait for Clk_period;
		Addr <=  "00000111011110";
		Trees_din <= x"006707a9";
		wait for Clk_period;
		Addr <=  "00000111011111";
		Trees_din <= x"01184308";
		wait for Clk_period;
		Addr <=  "00000111100000";
		Trees_din <= x"03029904";
		wait for Clk_period;
		Addr <=  "00000111100001";
		Trees_din <= x"007707a9";
		wait for Clk_period;
		Addr <=  "00000111100010";
		Trees_din <= x"ffb707a9";
		wait for Clk_period;
		Addr <=  "00000111100011";
		Trees_din <= x"0615fc04";
		wait for Clk_period;
		Addr <=  "00000111100100";
		Trees_din <= x"009507a9";
		wait for Clk_period;
		Addr <=  "00000111100101";
		Trees_din <= x"003007a9";
		wait for Clk_period;
		Addr <=  "00000111100110";
		Trees_din <= x"ff9a07a9";
		wait for Clk_period;
		Addr <=  "00000111100111";
		Trees_din <= x"03092d04";
		wait for Clk_period;
		Addr <=  "00000111101000";
		Trees_din <= x"ff9107a9";
		wait for Clk_period;
		Addr <=  "00000111101001";
		Trees_din <= x"000e07a9";
		wait for Clk_period;
		Addr <=  "00000111101010";
		Trees_din <= x"01096520";
		wait for Clk_period;
		Addr <=  "00000111101011";
		Trees_din <= x"10fc6f08";
		wait for Clk_period;
		Addr <=  "00000111101100";
		Trees_din <= x"1a005104";
		wait for Clk_period;
		Addr <=  "00000111101101";
		Trees_din <= x"ffa10825";
		wait for Clk_period;
		Addr <=  "00000111101110";
		Trees_din <= x"006d0825";
		wait for Clk_period;
		Addr <=  "00000111101111";
		Trees_din <= x"0105190c";
		wait for Clk_period;
		Addr <=  "00000111110000";
		Trees_din <= x"0ef83c08";
		wait for Clk_period;
		Addr <=  "00000111110001";
		Trees_din <= x"08005204";
		wait for Clk_period;
		Addr <=  "00000111110010";
		Trees_din <= x"00480825";
		wait for Clk_period;
		Addr <=  "00000111110011";
		Trees_din <= x"ffa20825";
		wait for Clk_period;
		Addr <=  "00000111110100";
		Trees_din <= x"ff680825";
		wait for Clk_period;
		Addr <=  "00000111110101";
		Trees_din <= x"00fdf108";
		wait for Clk_period;
		Addr <=  "00000111110110";
		Trees_din <= x"06fe4104";
		wait for Clk_period;
		Addr <=  "00000111110111";
		Trees_din <= x"fff00825";
		wait for Clk_period;
		Addr <=  "00000111111000";
		Trees_din <= x"ff920825";
		wait for Clk_period;
		Addr <=  "00000111111001";
		Trees_din <= x"00460825";
		wait for Clk_period;
		Addr <=  "00000111111010";
		Trees_din <= x"021cf41c";
		wait for Clk_period;
		Addr <=  "00000111111011";
		Trees_din <= x"061cb518";
		wait for Clk_period;
		Addr <=  "00000111111100";
		Trees_din <= x"01184310";
		wait for Clk_period;
		Addr <=  "00000111111101";
		Trees_din <= x"03010308";
		wait for Clk_period;
		Addr <=  "00000111111110";
		Trees_din <= x"05fb0d04";
		wait for Clk_period;
		Addr <=  "00000111111111";
		Trees_din <= x"fff20825";
		wait for Clk_period;
		Addr <=  "00001000000000";
		Trees_din <= x"006a0825";
		wait for Clk_period;
		Addr <=  "00001000000001";
		Trees_din <= x"0b020804";
		wait for Clk_period;
		Addr <=  "00001000000010";
		Trees_din <= x"ff940825";
		wait for Clk_period;
		Addr <=  "00001000000011";
		Trees_din <= x"001f0825";
		wait for Clk_period;
		Addr <=  "00001000000100";
		Trees_din <= x"1c002704";
		wait for Clk_period;
		Addr <=  "00001000000101";
		Trees_din <= x"00300825";
		wait for Clk_period;
		Addr <=  "00001000000110";
		Trees_din <= x"008f0825";
		wait for Clk_period;
		Addr <=  "00001000000111";
		Trees_din <= x"ffa30825";
		wait for Clk_period;
		Addr <=  "00001000001000";
		Trees_din <= x"ff9f0825";
		wait for Clk_period;
		Addr <=  "00001000001001";
		Trees_din <= x"010d0428";
		wait for Clk_period;
		Addr <=  "00001000001010";
		Trees_din <= x"01051914";
		wait for Clk_period;
		Addr <=  "00001000001011";
		Trees_din <= x"10fc6f08";
		wait for Clk_period;
		Addr <=  "00001000001100";
		Trees_din <= x"01fe1c04";
		wait for Clk_period;
		Addr <=  "00001000001101";
		Trees_din <= x"ffa908b1";
		wait for Clk_period;
		Addr <=  "00001000001110";
		Trees_din <= x"006608b1";
		wait for Clk_period;
		Addr <=  "00001000001111";
		Trees_din <= x"0ef83c08";
		wait for Clk_period;
		Addr <=  "00001000010000";
		Trees_din <= x"08005204";
		wait for Clk_period;
		Addr <=  "00001000010001";
		Trees_din <= x"004608b1";
		wait for Clk_period;
		Addr <=  "00001000010010";
		Trees_din <= x"ffaa08b1";
		wait for Clk_period;
		Addr <=  "00001000010011";
		Trees_din <= x"ff6908b1";
		wait for Clk_period;
		Addr <=  "00001000010100";
		Trees_din <= x"00f56608";
		wait for Clk_period;
		Addr <=  "00001000010101";
		Trees_din <= x"16031e04";
		wait for Clk_period;
		Addr <=  "00001000010110";
		Trees_din <= x"ff8608b1";
		wait for Clk_period;
		Addr <=  "00001000010111";
		Trees_din <= x"000008b1";
		wait for Clk_period;
		Addr <=  "00001000011000";
		Trees_din <= x"0c01b808";
		wait for Clk_period;
		Addr <=  "00001000011001";
		Trees_din <= x"08005304";
		wait for Clk_period;
		Addr <=  "00001000011010";
		Trees_din <= x"000908b1";
		wait for Clk_period;
		Addr <=  "00001000011011";
		Trees_din <= x"005f08b1";
		wait for Clk_period;
		Addr <=  "00001000011100";
		Trees_din <= x"ffc108b1";
		wait for Clk_period;
		Addr <=  "00001000011101";
		Trees_din <= x"021a0318";
		wait for Clk_period;
		Addr <=  "00001000011110";
		Trees_din <= x"0614d410";
		wait for Clk_period;
		Addr <=  "00001000011111";
		Trees_din <= x"04121008";
		wait for Clk_period;
		Addr <=  "00001000100000";
		Trees_din <= x"05098d04";
		wait for Clk_period;
		Addr <=  "00001000100001";
		Trees_din <= x"008208b1";
		wait for Clk_period;
		Addr <=  "00001000100010";
		Trees_din <= x"002408b1";
		wait for Clk_period;
		Addr <=  "00001000100011";
		Trees_din <= x"01184304";
		wait for Clk_period;
		Addr <=  "00001000100100";
		Trees_din <= x"ffa808b1";
		wait for Clk_period;
		Addr <=  "00001000100101";
		Trees_din <= x"005b08b1";
		wait for Clk_period;
		Addr <=  "00001000100110";
		Trees_din <= x"0123d704";
		wait for Clk_period;
		Addr <=  "00001000100111";
		Trees_din <= x"ffa008b1";
		wait for Clk_period;
		Addr <=  "00001000101000";
		Trees_din <= x"003a08b1";
		wait for Clk_period;
		Addr <=  "00001000101001";
		Trees_din <= x"18003e04";
		wait for Clk_period;
		Addr <=  "00001000101010";
		Trees_din <= x"ffa508b1";
		wait for Clk_period;
		Addr <=  "00001000101011";
		Trees_din <= x"001308b1";
		wait for Clk_period;
		Addr <=  "00001000101100";
		Trees_din <= x"01081b1c";
		wait for Clk_period;
		Addr <=  "00001000101101";
		Trees_din <= x"10fc6f08";
		wait for Clk_period;
		Addr <=  "00001000101110";
		Trees_din <= x"01fe1c04";
		wait for Clk_period;
		Addr <=  "00001000101111";
		Trees_din <= x"ffb10925";
		wait for Clk_period;
		Addr <=  "00001000110000";
		Trees_din <= x"00590925";
		wait for Clk_period;
		Addr <=  "00001000110001";
		Trees_din <= x"0ef83c08";
		wait for Clk_period;
		Addr <=  "00001000110010";
		Trees_din <= x"14033804";
		wait for Clk_period;
		Addr <=  "00001000110011";
		Trees_din <= x"00450925";
		wait for Clk_period;
		Addr <=  "00001000110100";
		Trees_din <= x"ffae0925";
		wait for Clk_period;
		Addr <=  "00001000110101";
		Trees_din <= x"01051904";
		wait for Clk_period;
		Addr <=  "00001000110110";
		Trees_din <= x"ff6a0925";
		wait for Clk_period;
		Addr <=  "00001000110111";
		Trees_din <= x"00f95f04";
		wait for Clk_period;
		Addr <=  "00001000111000";
		Trees_din <= x"ff9f0925";
		wait for Clk_period;
		Addr <=  "00001000111001";
		Trees_din <= x"001f0925";
		wait for Clk_period;
		Addr <=  "00001000111010";
		Trees_din <= x"0116f118";
		wait for Clk_period;
		Addr <=  "00001000111011";
		Trees_din <= x"04073410";
		wait for Clk_period;
		Addr <=  "00001000111100";
		Trees_din <= x"060af00c";
		wait for Clk_period;
		Addr <=  "00001000111101";
		Trees_din <= x"15f9bc04";
		wait for Clk_period;
		Addr <=  "00001000111110";
		Trees_din <= x"ffed0925";
		wait for Clk_period;
		Addr <=  "00001000111111";
		Trees_din <= x"020b1e04";
		wait for Clk_period;
		Addr <=  "00001001000000";
		Trees_din <= x"00730925";
		wait for Clk_period;
		Addr <=  "00001001000001";
		Trees_din <= x"000e0925";
		wait for Clk_period;
		Addr <=  "00001001000010";
		Trees_din <= x"ffd60925";
		wait for Clk_period;
		Addr <=  "00001001000011";
		Trees_din <= x"0b020d04";
		wait for Clk_period;
		Addr <=  "00001001000100";
		Trees_din <= x"ff940925";
		wait for Clk_period;
		Addr <=  "00001001000101";
		Trees_din <= x"ffe30925";
		wait for Clk_period;
		Addr <=  "00001001000110";
		Trees_din <= x"050fb304";
		wait for Clk_period;
		Addr <=  "00001001000111";
		Trees_din <= x"006e0925";
		wait for Clk_period;
		Addr <=  "00001001001000";
		Trees_din <= x"ffdc0925";
		wait for Clk_period;
		Addr <=  "00001001001001";
		Trees_din <= x"010d0420";
		wait for Clk_period;
		Addr <=  "00001001001010";
		Trees_din <= x"000bb81c";
		wait for Clk_period;
		Addr <=  "00001001001011";
		Trees_din <= x"11003908";
		wait for Clk_period;
		Addr <=  "00001001001100";
		Trees_din <= x"12008904";
		wait for Clk_period;
		Addr <=  "00001001001101";
		Trees_din <= x"007c0999";
		wait for Clk_period;
		Addr <=  "00001001001110";
		Trees_din <= x"ffb80999";
		wait for Clk_period;
		Addr <=  "00001001001111";
		Trees_din <= x"01051908";
		wait for Clk_period;
		Addr <=  "00001001010000";
		Trees_din <= x"1a005104";
		wait for Clk_period;
		Addr <=  "00001001010001";
		Trees_din <= x"ff790999";
		wait for Clk_period;
		Addr <=  "00001001010010";
		Trees_din <= x"ffec0999";
		wait for Clk_period;
		Addr <=  "00001001010011";
		Trees_din <= x"0c00ba08";
		wait for Clk_period;
		Addr <=  "00001001010100";
		Trees_din <= x"03fd6d04";
		wait for Clk_period;
		Addr <=  "00001001010101";
		Trees_din <= x"00420999";
		wait for Clk_period;
		Addr <=  "00001001010110";
		Trees_din <= x"ffcd0999";
		wait for Clk_period;
		Addr <=  "00001001010111";
		Trees_din <= x"ffa00999";
		wait for Clk_period;
		Addr <=  "00001001011000";
		Trees_din <= x"ff6e0999";
		wait for Clk_period;
		Addr <=  "00001001011001";
		Trees_din <= x"0615fc14";
		wait for Clk_period;
		Addr <=  "00001001011010";
		Trees_din <= x"02160e0c";
		wait for Clk_period;
		Addr <=  "00001001011011";
		Trees_din <= x"04121008";
		wait for Clk_period;
		Addr <=  "00001001011100";
		Trees_din <= x"0110ce04";
		wait for Clk_period;
		Addr <=  "00001001011101";
		Trees_din <= x"002f0999";
		wait for Clk_period;
		Addr <=  "00001001011110";
		Trees_din <= x"00800999";
		wait for Clk_period;
		Addr <=  "00001001011111";
		Trees_din <= x"fffe0999";
		wait for Clk_period;
		Addr <=  "00001001100000";
		Trees_din <= x"04121004";
		wait for Clk_period;
		Addr <=  "00001001100001";
		Trees_din <= x"ffb70999";
		wait for Clk_period;
		Addr <=  "00001001100010";
		Trees_din <= x"001d0999";
		wait for Clk_period;
		Addr <=  "00001001100011";
		Trees_din <= x"0413db04";
		wait for Clk_period;
		Addr <=  "00001001100100";
		Trees_din <= x"ffb00999";
		wait for Clk_period;
		Addr <=  "00001001100101";
		Trees_din <= x"000f0999";
		wait for Clk_period;
		Addr <=  "00001001100110";
		Trees_din <= x"01081b14";
		wait for Clk_period;
		Addr <=  "00001001100111";
		Trees_din <= x"10fc6f04";
		wait for Clk_period;
		Addr <=  "00001001101000";
		Trees_din <= x"001809fd";
		wait for Clk_period;
		Addr <=  "00001001101001";
		Trees_din <= x"0c03860c";
		wait for Clk_period;
		Addr <=  "00001001101010";
		Trees_din <= x"01051904";
		wait for Clk_period;
		Addr <=  "00001001101011";
		Trees_din <= x"ff6e09fd";
		wait for Clk_period;
		Addr <=  "00001001101100";
		Trees_din <= x"00f95f04";
		wait for Clk_period;
		Addr <=  "00001001101101";
		Trees_din <= x"ffac09fd";
		wait for Clk_period;
		Addr <=  "00001001101110";
		Trees_din <= x"001a09fd";
		wait for Clk_period;
		Addr <=  "00001001101111";
		Trees_din <= x"000a09fd";
		wait for Clk_period;
		Addr <=  "00001001110000";
		Trees_din <= x"01184314";
		wait for Clk_period;
		Addr <=  "00001001110001";
		Trees_din <= x"0407890c";
		wait for Clk_period;
		Addr <=  "00001001110010";
		Trees_din <= x"010d0408";
		wait for Clk_period;
		Addr <=  "00001001110011";
		Trees_din <= x"0efdf604";
		wait for Clk_period;
		Addr <=  "00001001110100";
		Trees_din <= x"003609fd";
		wait for Clk_period;
		Addr <=  "00001001110101";
		Trees_din <= x"ffc809fd";
		wait for Clk_period;
		Addr <=  "00001001110110";
		Trees_din <= x"005a09fd";
		wait for Clk_period;
		Addr <=  "00001001110111";
		Trees_din <= x"0b020804";
		wait for Clk_period;
		Addr <=  "00001001111000";
		Trees_din <= x"ff9e09fd";
		wait for Clk_period;
		Addr <=  "00001001111001";
		Trees_din <= x"000509fd";
		wait for Clk_period;
		Addr <=  "00001001111010";
		Trees_din <= x"00c00004";
		wait for Clk_period;
		Addr <=  "00001001111011";
		Trees_din <= x"001909fd";
		wait for Clk_period;
		Addr <=  "00001001111100";
		Trees_din <= x"1602f904";
		wait for Clk_period;
		Addr <=  "00001001111101";
		Trees_din <= x"007509fd";
		wait for Clk_period;
		Addr <=  "00001001111110";
		Trees_din <= x"002009fd";
		wait for Clk_period;
		Addr <=  "00001001111111";
		Trees_din <= x"01081b14";
		wait for Clk_period;
		Addr <=  "00001010000000";
		Trees_din <= x"10fc6f04";
		wait for Clk_period;
		Addr <=  "00001010000001";
		Trees_din <= x"00180a51";
		wait for Clk_period;
		Addr <=  "00001010000010";
		Trees_din <= x"0ef83c04";
		wait for Clk_period;
		Addr <=  "00001010000011";
		Trees_din <= x"00110a51";
		wait for Clk_period;
		Addr <=  "00001010000100";
		Trees_din <= x"01051904";
		wait for Clk_period;
		Addr <=  "00001010000101";
		Trees_din <= x"ff700a51";
		wait for Clk_period;
		Addr <=  "00001010000110";
		Trees_din <= x"15fb4404";
		wait for Clk_period;
		Addr <=  "00001010000111";
		Trees_din <= x"00120a51";
		wait for Clk_period;
		Addr <=  "00001010001000";
		Trees_din <= x"ffb90a51";
		wait for Clk_period;
		Addr <=  "00001010001001";
		Trees_din <= x"050fb314";
		wait for Clk_period;
		Addr <=  "00001010001010";
		Trees_din <= x"011fa010";
		wait for Clk_period;
		Addr <=  "00001010001011";
		Trees_din <= x"060f950c";
		wait for Clk_period;
		Addr <=  "00001010001100";
		Trees_din <= x"0211e908";
		wait for Clk_period;
		Addr <=  "00001010001101";
		Trees_din <= x"0c02f904";
		wait for Clk_period;
		Addr <=  "00001010001110";
		Trees_din <= x"005b0a51";
		wait for Clk_period;
		Addr <=  "00001010001111";
		Trees_din <= x"fffe0a51";
		wait for Clk_period;
		Addr <=  "00001010010000";
		Trees_din <= x"ffb30a51";
		wait for Clk_period;
		Addr <=  "00001010010001";
		Trees_din <= x"ffa10a51";
		wait for Clk_period;
		Addr <=  "00001010010010";
		Trees_din <= x"00770a51";
		wait for Clk_period;
		Addr <=  "00001010010011";
		Trees_din <= x"ffc50a51";
		wait for Clk_period;
		Addr <=  "00001010010100";
		Trees_din <= x"010db61c";
		wait for Clk_period;
		Addr <=  "00001010010101";
		Trees_din <= x"000bb818";
		wait for Clk_period;
		Addr <=  "00001010010110";
		Trees_din <= x"12008e0c";
		wait for Clk_period;
		Addr <=  "00001010010111";
		Trees_din <= x"00020804";
		wait for Clk_period;
		Addr <=  "00001010011000";
		Trees_din <= x"ffc10ab5";
		wait for Clk_period;
		Addr <=  "00001010011001";
		Trees_din <= x"09027a04";
		wait for Clk_period;
		Addr <=  "00001010011010";
		Trees_din <= x"007c0ab5";
		wait for Clk_period;
		Addr <=  "00001010011011";
		Trees_din <= x"00030ab5";
		wait for Clk_period;
		Addr <=  "00001010011100";
		Trees_din <= x"01096508";
		wait for Clk_period;
		Addr <=  "00001010011101";
		Trees_din <= x"16037304";
		wait for Clk_period;
		Addr <=  "00001010011110";
		Trees_din <= x"ff840ab5";
		wait for Clk_period;
		Addr <=  "00001010011111";
		Trees_din <= x"fff30ab5";
		wait for Clk_period;
		Addr <=  "00001010100000";
		Trees_din <= x"fffa0ab5";
		wait for Clk_period;
		Addr <=  "00001010100001";
		Trees_din <= x"ff770ab5";
		wait for Clk_period;
		Addr <=  "00001010100010";
		Trees_din <= x"050fb314";
		wait for Clk_period;
		Addr <=  "00001010100011";
		Trees_din <= x"0615fc10";
		wait for Clk_period;
		Addr <=  "00001010100100";
		Trees_din <= x"0118430c";
		wait for Clk_period;
		Addr <=  "00001010100101";
		Trees_din <= x"0407d104";
		wait for Clk_period;
		Addr <=  "00001010100110";
		Trees_din <= x"005f0ab5";
		wait for Clk_period;
		Addr <=  "00001010100111";
		Trees_din <= x"0b01d204";
		wait for Clk_period;
		Addr <=  "00001010101000";
		Trees_din <= x"ffc00ab5";
		wait for Clk_period;
		Addr <=  "00001010101001";
		Trees_din <= x"00020ab5";
		wait for Clk_period;
		Addr <=  "00001010101010";
		Trees_din <= x"00750ab5";
		wait for Clk_period;
		Addr <=  "00001010101011";
		Trees_din <= x"ffea0ab5";
		wait for Clk_period;
		Addr <=  "00001010101100";
		Trees_din <= x"ffd90ab5";
		wait for Clk_period;
		Addr <=  "00001010101101";
		Trees_din <= x"010db620";
		wait for Clk_period;
		Addr <=  "00001010101110";
		Trees_din <= x"000bb81c";
		wait for Clk_period;
		Addr <=  "00001010101111";
		Trees_din <= x"11003908";
		wait for Clk_period;
		Addr <=  "00001010110000";
		Trees_din <= x"06fe4104";
		wait for Clk_period;
		Addr <=  "00001010110001";
		Trees_din <= x"004d0b19";
		wait for Clk_period;
		Addr <=  "00001010110010";
		Trees_din <= x"fff70b19";
		wait for Clk_period;
		Addr <=  "00001010110011";
		Trees_din <= x"01051908";
		wait for Clk_period;
		Addr <=  "00001010110100";
		Trees_din <= x"1a004f04";
		wait for Clk_period;
		Addr <=  "00001010110101";
		Trees_din <= x"ff8c0b19";
		wait for Clk_period;
		Addr <=  "00001010110110";
		Trees_din <= x"fff10b19";
		wait for Clk_period;
		Addr <=  "00001010110111";
		Trees_din <= x"00e9ab04";
		wait for Clk_period;
		Addr <=  "00001010111000";
		Trees_din <= x"ffad0b19";
		wait for Clk_period;
		Addr <=  "00001010111001";
		Trees_din <= x"0c00ba04";
		wait for Clk_period;
		Addr <=  "00001010111010";
		Trees_din <= x"00350b19";
		wait for Clk_period;
		Addr <=  "00001010111011";
		Trees_din <= x"ffd10b19";
		wait for Clk_period;
		Addr <=  "00001010111100";
		Trees_din <= x"ff7b0b19";
		wait for Clk_period;
		Addr <=  "00001010111101";
		Trees_din <= x"040ebb08";
		wait for Clk_period;
		Addr <=  "00001010111110";
		Trees_din <= x"0302e404";
		wait for Clk_period;
		Addr <=  "00001010111111";
		Trees_din <= x"005f0b19";
		wait for Clk_period;
		Addr <=  "00001011000000";
		Trees_din <= x"00050b19";
		wait for Clk_period;
		Addr <=  "00001011000001";
		Trees_din <= x"011fa004";
		wait for Clk_period;
		Addr <=  "00001011000010";
		Trees_din <= x"ffae0b19";
		wait for Clk_period;
		Addr <=  "00001011000011";
		Trees_din <= x"1402a104";
		wait for Clk_period;
		Addr <=  "00001011000100";
		Trees_din <= x"00110b19";
		wait for Clk_period;
		Addr <=  "00001011000101";
		Trees_din <= x"005c0b19";
		wait for Clk_period;
		Addr <=  "00001011000110";
		Trees_din <= x"010d0414";
		wait for Clk_period;
		Addr <=  "00001011000111";
		Trees_din <= x"10fc6f04";
		wait for Clk_period;
		Addr <=  "00001011001000";
		Trees_din <= x"001e0b65";
		wait for Clk_period;
		Addr <=  "00001011001001";
		Trees_din <= x"0ef85404";
		wait for Clk_period;
		Addr <=  "00001011001010";
		Trees_din <= x"00170b65";
		wait for Clk_period;
		Addr <=  "00001011001011";
		Trees_din <= x"01051904";
		wait for Clk_period;
		Addr <=  "00001011001100";
		Trees_din <= x"ff780b65";
		wait for Clk_period;
		Addr <=  "00001011001101";
		Trees_din <= x"0c00ba04";
		wait for Clk_period;
		Addr <=  "00001011001110";
		Trees_din <= x"00120b65";
		wait for Clk_period;
		Addr <=  "00001011001111";
		Trees_din <= x"ffb70b65";
		wait for Clk_period;
		Addr <=  "00001011010000";
		Trees_din <= x"0116f108";
		wait for Clk_period;
		Addr <=  "00001011010001";
		Trees_din <= x"0407d104";
		wait for Clk_period;
		Addr <=  "00001011010010";
		Trees_din <= x"00430b65";
		wait for Clk_period;
		Addr <=  "00001011010011";
		Trees_din <= x"ffba0b65";
		wait for Clk_period;
		Addr <=  "00001011010100";
		Trees_din <= x"09054708";
		wait for Clk_period;
		Addr <=  "00001011010101";
		Trees_din <= x"011fa004";
		wait for Clk_period;
		Addr <=  "00001011010110";
		Trees_din <= x"00230b65";
		wait for Clk_period;
		Addr <=  "00001011010111";
		Trees_din <= x"00670b65";
		wait for Clk_period;
		Addr <=  "00001011011000";
		Trees_din <= x"000a0b65";
		wait for Clk_period;
		Addr <=  "00001011011001";
		Trees_din <= x"0112461c";
		wait for Clk_period;
		Addr <=  "00001011011010";
		Trees_din <= x"03fdbf10";
		wait for Clk_period;
		Addr <=  "00001011011011";
		Trees_din <= x"12008e08";
		wait for Clk_period;
		Addr <=  "00001011011100";
		Trees_din <= x"11003904";
		wait for Clk_period;
		Addr <=  "00001011011101";
		Trees_din <= x"00590bb9";
		wait for Clk_period;
		Addr <=  "00001011011110";
		Trees_din <= x"fff00bb9";
		wait for Clk_period;
		Addr <=  "00001011011111";
		Trees_din <= x"01096504";
		wait for Clk_period;
		Addr <=  "00001011100000";
		Trees_din <= x"ffa00bb9";
		wait for Clk_period;
		Addr <=  "00001011100001";
		Trees_din <= x"002b0bb9";
		wait for Clk_period;
		Addr <=  "00001011100010";
		Trees_din <= x"01069b04";
		wait for Clk_period;
		Addr <=  "00001011100011";
		Trees_din <= x"ff830bb9";
		wait for Clk_period;
		Addr <=  "00001011100100";
		Trees_din <= x"10021e04";
		wait for Clk_period;
		Addr <=  "00001011100101";
		Trees_din <= x"ffc10bb9";
		wait for Clk_period;
		Addr <=  "00001011100110";
		Trees_din <= x"00020bb9";
		wait for Clk_period;
		Addr <=  "00001011100111";
		Trees_din <= x"0410ae08";
		wait for Clk_period;
		Addr <=  "00001011101000";
		Trees_din <= x"0302e404";
		wait for Clk_period;
		Addr <=  "00001011101001";
		Trees_din <= x"00610bb9";
		wait for Clk_period;
		Addr <=  "00001011101010";
		Trees_din <= x"00110bb9";
		wait for Clk_period;
		Addr <=  "00001011101011";
		Trees_din <= x"16006c04";
		wait for Clk_period;
		Addr <=  "00001011101100";
		Trees_din <= x"ffdb0bb9";
		wait for Clk_period;
		Addr <=  "00001011101101";
		Trees_din <= x"003a0bb9";
		wait for Clk_period;
		Addr <=  "00001011101110";
		Trees_din <= x"010e9018";
		wait for Clk_period;
		Addr <=  "00001011101111";
		Trees_din <= x"03fdbf10";
		wait for Clk_period;
		Addr <=  "00001011110000";
		Trees_din <= x"0c02d60c";
		wait for Clk_period;
		Addr <=  "00001011110001";
		Trees_din <= x"01002704";
		wait for Clk_period;
		Addr <=  "00001011110010";
		Trees_din <= x"ff9c0c05";
		wait for Clk_period;
		Addr <=  "00001011110011";
		Trees_din <= x"19009204";
		wait for Clk_period;
		Addr <=  "00001011110100";
		Trees_din <= x"00260c05";
		wait for Clk_period;
		Addr <=  "00001011110101";
		Trees_din <= x"ffdd0c05";
		wait for Clk_period;
		Addr <=  "00001011110110";
		Trees_din <= x"00340c05";
		wait for Clk_period;
		Addr <=  "00001011110111";
		Trees_din <= x"02047404";
		wait for Clk_period;
		Addr <=  "00001011111000";
		Trees_din <= x"ff890c05";
		wait for Clk_period;
		Addr <=  "00001011111001";
		Trees_din <= x"ffda0c05";
		wait for Clk_period;
		Addr <=  "00001011111010";
		Trees_din <= x"040ebb08";
		wait for Clk_period;
		Addr <=  "00001011111011";
		Trees_din <= x"0302e404";
		wait for Clk_period;
		Addr <=  "00001011111100";
		Trees_din <= x"00530c05";
		wait for Clk_period;
		Addr <=  "00001011111101";
		Trees_din <= x"00090c05";
		wait for Clk_period;
		Addr <=  "00001011111110";
		Trees_din <= x"011fa004";
		wait for Clk_period;
		Addr <=  "00001011111111";
		Trees_din <= x"ffb90c05";
		wait for Clk_period;
		Addr <=  "00001100000000";
		Trees_din <= x"00420c05";
		wait for Clk_period;
		Addr <=  "00001100000001";
		Trees_din <= x"0112461c";
		wait for Clk_period;
		Addr <=  "00001100000010";
		Trees_din <= x"03fdbf10";
		wait for Clk_period;
		Addr <=  "00001100000011";
		Trees_din <= x"12008e08";
		wait for Clk_period;
		Addr <=  "00001100000100";
		Trees_din <= x"09027a04";
		wait for Clk_period;
		Addr <=  "00001100000101";
		Trees_din <= x"00490c51";
		wait for Clk_period;
		Addr <=  "00001100000110";
		Trees_din <= x"ffeb0c51";
		wait for Clk_period;
		Addr <=  "00001100000111";
		Trees_din <= x"01037504";
		wait for Clk_period;
		Addr <=  "00001100001000";
		Trees_din <= x"ffa30c51";
		wait for Clk_period;
		Addr <=  "00001100001001";
		Trees_din <= x"00050c51";
		wait for Clk_period;
		Addr <=  "00001100001010";
		Trees_din <= x"01069b04";
		wait for Clk_period;
		Addr <=  "00001100001011";
		Trees_din <= x"ff8e0c51";
		wait for Clk_period;
		Addr <=  "00001100001100";
		Trees_din <= x"0d019f04";
		wait for Clk_period;
		Addr <=  "00001100001101";
		Trees_din <= x"fffa0c51";
		wait for Clk_period;
		Addr <=  "00001100001110";
		Trees_din <= x"ffd00c51";
		wait for Clk_period;
		Addr <=  "00001100001111";
		Trees_din <= x"040ebb04";
		wait for Clk_period;
		Addr <=  "00001100010000";
		Trees_din <= x"004a0c51";
		wait for Clk_period;
		Addr <=  "00001100010001";
		Trees_din <= x"16006c04";
		wait for Clk_period;
		Addr <=  "00001100010010";
		Trees_din <= x"ffeb0c51";
		wait for Clk_period;
		Addr <=  "00001100010011";
		Trees_din <= x"002e0c51";
		wait for Clk_period;
		Addr <=  "00001100010100";
		Trees_din <= x"01124618";
		wait for Clk_period;
		Addr <=  "00001100010101";
		Trees_din <= x"03fdbf10";
		wait for Clk_period;
		Addr <=  "00001100010110";
		Trees_din <= x"12008e08";
		wait for Clk_period;
		Addr <=  "00001100010111";
		Trees_din <= x"1e007704";
		wait for Clk_period;
		Addr <=  "00001100011000";
		Trees_din <= x"00430c95";
		wait for Clk_period;
		Addr <=  "00001100011001";
		Trees_din <= x"fff50c95";
		wait for Clk_period;
		Addr <=  "00001100011010";
		Trees_din <= x"01037504";
		wait for Clk_period;
		Addr <=  "00001100011011";
		Trees_din <= x"ffa90c95";
		wait for Clk_period;
		Addr <=  "00001100011100";
		Trees_din <= x"00050c95";
		wait for Clk_period;
		Addr <=  "00001100011101";
		Trees_din <= x"01069b04";
		wait for Clk_period;
		Addr <=  "00001100011110";
		Trees_din <= x"ff940c95";
		wait for Clk_period;
		Addr <=  "00001100011111";
		Trees_din <= x"ffdd0c95";
		wait for Clk_period;
		Addr <=  "00001100100000";
		Trees_din <= x"17004b08";
		wait for Clk_period;
		Addr <=  "00001100100001";
		Trees_din <= x"011cba04";
		wait for Clk_period;
		Addr <=  "00001100100010";
		Trees_din <= x"000d0c95";
		wait for Clk_period;
		Addr <=  "00001100100011";
		Trees_din <= x"00560c95";
		wait for Clk_period;
		Addr <=  "00001100100100";
		Trees_din <= x"ffff0c95";
		wait for Clk_period;
		Addr <=  "00001100100101";
		Trees_din <= x"01124618";
		wait for Clk_period;
		Addr <=  "00001100100110";
		Trees_din <= x"11008308";
		wait for Clk_period;
		Addr <=  "00001100100111";
		Trees_din <= x"11003604";
		wait for Clk_period;
		Addr <=  "00001100101000";
		Trees_din <= x"ffc60cd9";
		wait for Clk_period;
		Addr <=  "00001100101001";
		Trees_din <= x"00340cd9";
		wait for Clk_period;
		Addr <=  "00001100101010";
		Trees_din <= x"03fcb608";
		wait for Clk_period;
		Addr <=  "00001100101011";
		Trees_din <= x"0f00f504";
		wait for Clk_period;
		Addr <=  "00001100101100";
		Trees_din <= x"00170cd9";
		wait for Clk_period;
		Addr <=  "00001100101101";
		Trees_din <= x"ffd10cd9";
		wait for Clk_period;
		Addr <=  "00001100101110";
		Trees_din <= x"1403a604";
		wait for Clk_period;
		Addr <=  "00001100101111";
		Trees_din <= x"ff980cd9";
		wait for Clk_period;
		Addr <=  "00001100110000";
		Trees_din <= x"ffe20cd9";
		wait for Clk_period;
		Addr <=  "00001100110001";
		Trees_din <= x"011fa008";
		wait for Clk_period;
		Addr <=  "00001100110010";
		Trees_din <= x"00c00004";
		wait for Clk_period;
		Addr <=  "00001100110011";
		Trees_din <= x"ffd10cd9";
		wait for Clk_period;
		Addr <=  "00001100110100";
		Trees_din <= x"003e0cd9";
		wait for Clk_period;
		Addr <=  "00001100110101";
		Trees_din <= x"00480cd9";
		wait for Clk_period;
		Addr <=  "00001100110110";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00001100110111";
		Trees_din <= x"010d0410";
		wait for Clk_period;
		Addr <=  "00001100111000";
		Trees_din <= x"11003904";
		wait for Clk_period;
		Addr <=  "00001100111001";
		Trees_din <= x"000f0d19";
		wait for Clk_period;
		Addr <=  "00001100111010";
		Trees_din <= x"01051904";
		wait for Clk_period;
		Addr <=  "00001100111011";
		Trees_din <= x"ff9f0d19";
		wait for Clk_period;
		Addr <=  "00001100111100";
		Trees_din <= x"14032d04";
		wait for Clk_period;
		Addr <=  "00001100111101";
		Trees_din <= x"ffd10d19";
		wait for Clk_period;
		Addr <=  "00001100111110";
		Trees_din <= x"00180d19";
		wait for Clk_period;
		Addr <=  "00001100111111";
		Trees_din <= x"01184308";
		wait for Clk_period;
		Addr <=  "00001101000000";
		Trees_din <= x"0407d104";
		wait for Clk_period;
		Addr <=  "00001101000001";
		Trees_din <= x"00370d19";
		wait for Clk_period;
		Addr <=  "00001101000010";
		Trees_din <= x"ffd20d19";
		wait for Clk_period;
		Addr <=  "00001101000011";
		Trees_din <= x"00c00004";
		wait for Clk_period;
		Addr <=  "00001101000100";
		Trees_din <= x"000c0d19";
		wait for Clk_period;
		Addr <=  "00001101000101";
		Trees_din <= x"00490d19";
		wait for Clk_period;
		Addr <=  "00001101000110";
		Trees_din <= x"010d0410";
		wait for Clk_period;
		Addr <=  "00001101000111";
		Trees_din <= x"12008e08";
		wait for Clk_period;
		Addr <=  "00001101001000";
		Trees_din <= x"18003e04";
		wait for Clk_period;
		Addr <=  "00001101001001";
		Trees_din <= x"00310d55";
		wait for Clk_period;
		Addr <=  "00001101001010";
		Trees_din <= x"ffdd0d55";
		wait for Clk_period;
		Addr <=  "00001101001011";
		Trees_din <= x"01069b04";
		wait for Clk_period;
		Addr <=  "00001101001100";
		Trees_din <= x"ff9d0d55";
		wait for Clk_period;
		Addr <=  "00001101001101";
		Trees_din <= x"fff50d55";
		wait for Clk_period;
		Addr <=  "00001101001110";
		Trees_din <= x"011fa00c";
		wait for Clk_period;
		Addr <=  "00001101001111";
		Trees_din <= x"040db708";
		wait for Clk_period;
		Addr <=  "00001101010000";
		Trees_din <= x"03005904";
		wait for Clk_period;
		Addr <=  "00001101010001";
		Trees_din <= x"003f0d55";
		wait for Clk_period;
		Addr <=  "00001101010010";
		Trees_din <= x"00070d55";
		wait for Clk_period;
		Addr <=  "00001101010011";
		Trees_din <= x"ffc50d55";
		wait for Clk_period;
		Addr <=  "00001101010100";
		Trees_din <= x"00420d55";
		wait for Clk_period;
		Addr <=  "00001101010101";
		Trees_din <= x"01124610";
		wait for Clk_period;
		Addr <=  "00001101010110";
		Trees_din <= x"03fdbf0c";
		wait for Clk_period;
		Addr <=  "00001101010111";
		Trees_din <= x"19009508";
		wait for Clk_period;
		Addr <=  "00001101011000";
		Trees_din <= x"18003e04";
		wait for Clk_period;
		Addr <=  "00001101011001";
		Trees_din <= x"00380d81";
		wait for Clk_period;
		Addr <=  "00001101011010";
		Trees_din <= x"fff20d81";
		wait for Clk_period;
		Addr <=  "00001101011011";
		Trees_din <= x"ffd30d81";
		wait for Clk_period;
		Addr <=  "00001101011100";
		Trees_din <= x"ffb80d81";
		wait for Clk_period;
		Addr <=  "00001101011101";
		Trees_din <= x"0fff0604";
		wait for Clk_period;
		Addr <=  "00001101011110";
		Trees_din <= x"00040d81";
		wait for Clk_period;
		Addr <=  "00001101011111";
		Trees_din <= x"00380d81";
		wait for Clk_period;
		Addr <=  "00001101100000";
		Trees_din <= x"010d0410";
		wait for Clk_period;
		Addr <=  "00001101100001";
		Trees_din <= x"12008e08";
		wait for Clk_period;
		Addr <=  "00001101100010";
		Trees_din <= x"09027a04";
		wait for Clk_period;
		Addr <=  "00001101100011";
		Trees_din <= x"00240db5";
		wait for Clk_period;
		Addr <=  "00001101100100";
		Trees_din <= x"ffe20db5";
		wait for Clk_period;
		Addr <=  "00001101100101";
		Trees_din <= x"01069b04";
		wait for Clk_period;
		Addr <=  "00001101100110";
		Trees_din <= x"ffa40db5";
		wait for Clk_period;
		Addr <=  "00001101100111";
		Trees_din <= x"fff90db5";
		wait for Clk_period;
		Addr <=  "00001101101000";
		Trees_din <= x"011fa008";
		wait for Clk_period;
		Addr <=  "00001101101001";
		Trees_din <= x"00c9cc04";
		wait for Clk_period;
		Addr <=  "00001101101010";
		Trees_din <= x"ffd90db5";
		wait for Clk_period;
		Addr <=  "00001101101011";
		Trees_din <= x"00340db5";
		wait for Clk_period;
		Addr <=  "00001101101100";
		Trees_din <= x"003d0db5";
		wait for Clk_period;
		Addr <=  "00001101101101";
		Trees_din <= x"01124610";
		wait for Clk_period;
		Addr <=  "00001101101110";
		Trees_din <= x"11008308";
		wait for Clk_period;
		Addr <=  "00001101101111";
		Trees_din <= x"09027b04";
		wait for Clk_period;
		Addr <=  "00001101110000";
		Trees_din <= x"00260de1";
		wait for Clk_period;
		Addr <=  "00001101110001";
		Trees_din <= x"ffe70de1";
		wait for Clk_period;
		Addr <=  "00001101110010";
		Trees_din <= x"03fcb604";
		wait for Clk_period;
		Addr <=  "00001101110011";
		Trees_din <= x"fff60de1";
		wait for Clk_period;
		Addr <=  "00001101110100";
		Trees_din <= x"ffb50de1";
		wait for Clk_period;
		Addr <=  "00001101110101";
		Trees_din <= x"01184304";
		wait for Clk_period;
		Addr <=  "00001101110110";
		Trees_din <= x"00050de1";
		wait for Clk_period;
		Addr <=  "00001101110111";
		Trees_din <= x"00350de1";
		wait for Clk_period;
		Addr <=  "00001101111000";
		Trees_din <= x"010d040c";
		wait for Clk_period;
		Addr <=  "00001101111001";
		Trees_din <= x"11003904";
		wait for Clk_period;
		Addr <=  "00001101111010";
		Trees_din <= x"000f0e0d";
		wait for Clk_period;
		Addr <=  "00001101111011";
		Trees_din <= x"01051904";
		wait for Clk_period;
		Addr <=  "00001101111100";
		Trees_din <= x"ffb20e0d";
		wait for Clk_period;
		Addr <=  "00001101111101";
		Trees_din <= x"fff70e0d";
		wait for Clk_period;
		Addr <=  "00001101111110";
		Trees_din <= x"040ebb08";
		wait for Clk_period;
		Addr <=  "00001101111111";
		Trees_din <= x"0a015d04";
		wait for Clk_period;
		Addr <=  "00001110000000";
		Trees_din <= x"003d0e0d";
		wait for Clk_period;
		Addr <=  "00001110000001";
		Trees_din <= x"00100e0d";
		wait for Clk_period;
		Addr <=  "00001110000010";
		Trees_din <= x"00000e0d";
		wait for Clk_period;
		Addr <=  "00001110000011";
		Trees_din <= x"01184310";
		wait for Clk_period;
		Addr <=  "00001110000100";
		Trees_din <= x"03ff770c";
		wait for Clk_period;
		Addr <=  "00001110000101";
		Trees_din <= x"01096508";
		wait for Clk_period;
		Addr <=  "00001110000110";
		Trees_din <= x"12008e04";
		wait for Clk_period;
		Addr <=  "00001110000111";
		Trees_din <= x"00130e31";
		wait for Clk_period;
		Addr <=  "00001110001000";
		Trees_din <= x"ffc10e31";
		wait for Clk_period;
		Addr <=  "00001110001001";
		Trees_din <= x"00280e31";
		wait for Clk_period;
		Addr <=  "00001110001010";
		Trees_din <= x"ffbf0e31";
		wait for Clk_period;
		Addr <=  "00001110001011";
		Trees_din <= x"00330e31";
		wait for Clk_period;
		Addr <=  "00001110001100";
		Trees_din <= x"0116f110";
		wait for Clk_period;
		Addr <=  "00001110001101";
		Trees_din <= x"03ff770c";
		wait for Clk_period;
		Addr <=  "00001110001110";
		Trees_din <= x"01096508";
		wait for Clk_period;
		Addr <=  "00001110001111";
		Trees_din <= x"12008e04";
		wait for Clk_period;
		Addr <=  "00001110010000";
		Trees_din <= x"00100e5d";
		wait for Clk_period;
		Addr <=  "00001110010001";
		Trees_din <= x"ffc60e5d";
		wait for Clk_period;
		Addr <=  "00001110010010";
		Trees_din <= x"00200e5d";
		wait for Clk_period;
		Addr <=  "00001110010011";
		Trees_din <= x"ffc00e5d";
		wait for Clk_period;
		Addr <=  "00001110010100";
		Trees_din <= x"011fa004";
		wait for Clk_period;
		Addr <=  "00001110010101";
		Trees_din <= x"000c0e5d";
		wait for Clk_period;
		Addr <=  "00001110010110";
		Trees_din <= x"00360e5d";
		wait for Clk_period;
		Addr <=  "00001110010111";
		Trees_din <= x"0112460c";
		wait for Clk_period;
		Addr <=  "00001110011000";
		Trees_din <= x"11008304";
		wait for Clk_period;
		Addr <=  "00001110011001";
		Trees_din <= x"00090e81";
		wait for Clk_period;
		Addr <=  "00001110011010";
		Trees_din <= x"03fcb604";
		wait for Clk_period;
		Addr <=  "00001110011011";
		Trees_din <= x"fff80e81";
		wait for Clk_period;
		Addr <=  "00001110011100";
		Trees_din <= x"ffbf0e81";
		wait for Clk_period;
		Addr <=  "00001110011101";
		Trees_din <= x"1401c704";
		wait for Clk_period;
		Addr <=  "00001110011110";
		Trees_din <= x"00060e81";
		wait for Clk_period;
		Addr <=  "00001110011111";
		Trees_din <= x"00320e81";
		wait for Clk_period;
		Addr <=  "00001110100000";
		Trees_din <= x"01184310";
		wait for Clk_period;
		Addr <=  "00001110100001";
		Trees_din <= x"03ff770c";
		wait for Clk_period;
		Addr <=  "00001110100010";
		Trees_din <= x"01096508";
		wait for Clk_period;
		Addr <=  "00001110100011";
		Trees_din <= x"12008e04";
		wait for Clk_period;
		Addr <=  "00001110100100";
		Trees_din <= x"000e0ea5";
		wait for Clk_period;
		Addr <=  "00001110100101";
		Trees_din <= x"ffcb0ea5";
		wait for Clk_period;
		Addr <=  "00001110100110";
		Trees_din <= x"00210ea5";
		wait for Clk_period;
		Addr <=  "00001110100111";
		Trees_din <= x"ffc80ea5";
		wait for Clk_period;
		Addr <=  "00001110101000";
		Trees_din <= x"002d0ea5";
		wait for Clk_period;
		Addr <=  "00001110101001";
		Trees_din <= x"010e900c";
		wait for Clk_period;
		Addr <=  "00001110101010";
		Trees_din <= x"11008304";
		wait for Clk_period;
		Addr <=  "00001110101011";
		Trees_din <= x"00060ec9";
		wait for Clk_period;
		Addr <=  "00001110101100";
		Trees_din <= x"0a00b004";
		wait for Clk_period;
		Addr <=  "00001110101101";
		Trees_din <= x"fff40ec9";
		wait for Clk_period;
		Addr <=  "00001110101110";
		Trees_din <= x"ffc50ec9";
		wait for Clk_period;
		Addr <=  "00001110101111";
		Trees_din <= x"040ebb04";
		wait for Clk_period;
		Addr <=  "00001110110000";
		Trees_din <= x"002f0ec9";
		wait for Clk_period;
		Addr <=  "00001110110001";
		Trees_din <= x"00020ec9";
		wait for Clk_period;
		Addr <=  "00001110110010";
		Trees_din <= x"01184310";
		wait for Clk_period;
		Addr <=  "00001110110011";
		Trees_din <= x"03ff770c";
		wait for Clk_period;
		Addr <=  "00001110110100";
		Trees_din <= x"01069b08";
		wait for Clk_period;
		Addr <=  "00001110110101";
		Trees_din <= x"09027a04";
		wait for Clk_period;
		Addr <=  "00001110110110";
		Trees_din <= x"00070eed";
		wait for Clk_period;
		Addr <=  "00001110110111";
		Trees_din <= x"ffd40eed";
		wait for Clk_period;
		Addr <=  "00001110111000";
		Trees_din <= x"001a0eed";
		wait for Clk_period;
		Addr <=  "00001110111001";
		Trees_din <= x"ffcc0eed";
		wait for Clk_period;
		Addr <=  "00001110111010";
		Trees_din <= x"002a0eed";
		wait for Clk_period;
		Addr <=  "00001110111011";
		Trees_din <= x"0112460c";
		wait for Clk_period;
		Addr <=  "00001110111100";
		Trees_din <= x"06ffd708";
		wait for Clk_period;
		Addr <=  "00001110111101";
		Trees_din <= x"06fe1a04";
		wait for Clk_period;
		Addr <=  "00001110111110";
		Trees_din <= x"ffec0f11";
		wait for Clk_period;
		Addr <=  "00001110111111";
		Trees_din <= x"00170f11";
		wait for Clk_period;
		Addr <=  "00001111000000";
		Trees_din <= x"ffd20f11";
		wait for Clk_period;
		Addr <=  "00001111000001";
		Trees_din <= x"011fa004";
		wait for Clk_period;
		Addr <=  "00001111000010";
		Trees_din <= x"00080f11";
		wait for Clk_period;
		Addr <=  "00001111000011";
		Trees_din <= x"00310f11";
		wait for Clk_period;
		Addr <=  "00001111000100";
		Trees_din <= x"010e900c";
		wait for Clk_period;
		Addr <=  "00001111000101";
		Trees_din <= x"11008304";
		wait for Clk_period;
		Addr <=  "00001111000110";
		Trees_din <= x"00040f35";
		wait for Clk_period;
		Addr <=  "00001111000111";
		Trees_din <= x"01037504";
		wait for Clk_period;
		Addr <=  "00001111001000";
		Trees_din <= x"ffcb0f35";
		wait for Clk_period;
		Addr <=  "00001111001001";
		Trees_din <= x"fff40f35";
		wait for Clk_period;
		Addr <=  "00001111001010";
		Trees_din <= x"16007104";
		wait for Clk_period;
		Addr <=  "00001111001011";
		Trees_din <= x"00030f35";
		wait for Clk_period;
		Addr <=  "00001111001100";
		Trees_din <= x"002f0f35";
		wait for Clk_period;
		Addr <=  "00001111001101";
		Trees_din <= x"0116f10c";
		wait for Clk_period;
		Addr <=  "00001111001110";
		Trees_din <= x"1101bb08";
		wait for Clk_period;
		Addr <=  "00001111001111";
		Trees_din <= x"19009904";
		wait for Clk_period;
		Addr <=  "00001111010000";
		Trees_din <= x"00180f59";
		wait for Clk_period;
		Addr <=  "00001111010001";
		Trees_din <= x"ffe40f59";
		wait for Clk_period;
		Addr <=  "00001111010010";
		Trees_din <= x"ffd40f59";
		wait for Clk_period;
		Addr <=  "00001111010011";
		Trees_din <= x"011fa004";
		wait for Clk_period;
		Addr <=  "00001111010100";
		Trees_din <= x"00070f59";
		wait for Clk_period;
		Addr <=  "00001111010101";
		Trees_din <= x"002f0f59";
		wait for Clk_period;
		Addr <=  "00001111010110";
		Trees_din <= x"010e9008";
		wait for Clk_period;
		Addr <=  "00001111010111";
		Trees_din <= x"06ffd004";
		wait for Clk_period;
		Addr <=  "00001111011000";
		Trees_din <= x"ffff0f75";
		wait for Clk_period;
		Addr <=  "00001111011001";
		Trees_din <= x"ffd20f75";
		wait for Clk_period;
		Addr <=  "00001111011010";
		Trees_din <= x"040ebb04";
		wait for Clk_period;
		Addr <=  "00001111011011";
		Trees_din <= x"002c0f75";
		wait for Clk_period;
		Addr <=  "00001111011100";
		Trees_din <= x"00010f75";
		wait for Clk_period;
		Addr <=  "00001111011101";
		Trees_din <= x"011a8c0c";
		wait for Clk_period;
		Addr <=  "00001111011110";
		Trees_din <= x"03fdbf08";
		wait for Clk_period;
		Addr <=  "00001111011111";
		Trees_din <= x"19009504";
		wait for Clk_period;
		Addr <=  "00001111100000";
		Trees_din <= x"00190f91";
		wait for Clk_period;
		Addr <=  "00001111100001";
		Trees_din <= x"ffeb0f91";
		wait for Clk_period;
		Addr <=  "00001111100010";
		Trees_din <= x"ffd90f91";
		wait for Clk_period;
		Addr <=  "00001111100011";
		Trees_din <= x"00280f91";
		wait for Clk_period;
		Addr <=  "00001111100100";
		Trees_din <= x"01069b04";
		wait for Clk_period;
		Addr <=  "00001111100101";
		Trees_din <= x"ffdd0fad";
		wait for Clk_period;
		Addr <=  "00001111100110";
		Trees_din <= x"07005404";
		wait for Clk_period;
		Addr <=  "00001111100111";
		Trees_din <= x"fff40fad";
		wait for Clk_period;
		Addr <=  "00001111101000";
		Trees_din <= x"1b025704";
		wait for Clk_period;
		Addr <=  "00001111101001";
		Trees_din <= x"00300fad";
		wait for Clk_period;
		Addr <=  "00001111101010";
		Trees_din <= x"ffff0fad";
		wait for Clk_period;
		Addr <=  "00001111101011";
		Trees_din <= x"01124608";
		wait for Clk_period;
		Addr <=  "00001111101100";
		Trees_din <= x"06ffd704";
		wait for Clk_period;
		Addr <=  "00001111101101";
		Trees_din <= x"00020fc9";
		wait for Clk_period;
		Addr <=  "00001111101110";
		Trees_din <= x"ffd80fc9";
		wait for Clk_period;
		Addr <=  "00001111101111";
		Trees_din <= x"011fa004";
		wait for Clk_period;
		Addr <=  "00001111110000";
		Trees_din <= x"00070fc9";
		wait for Clk_period;
		Addr <=  "00001111110001";
		Trees_din <= x"002d0fc9";
		wait for Clk_period;
		Addr <=  "00001111110010";
		Trees_din <= x"010d0408";
		wait for Clk_period;
		Addr <=  "00001111110011";
		Trees_din <= x"12008e04";
		wait for Clk_period;
		Addr <=  "00001111110100";
		Trees_din <= x"00050fe5";
		wait for Clk_period;
		Addr <=  "00001111110101";
		Trees_din <= x"ffd50fe5";
		wait for Clk_period;
		Addr <=  "00001111110110";
		Trees_din <= x"040ebb04";
		wait for Clk_period;
		Addr <=  "00001111110111";
		Trees_din <= x"00290fe5";
		wait for Clk_period;
		Addr <=  "00001111111000";
		Trees_din <= x"ffff0fe5";
		wait for Clk_period;
		Addr <=  "00001111111001";
		Trees_din <= x"01051904";
		wait for Clk_period;
		Addr <=  "00001111111010";
		Trees_din <= x"ffdd1001";
		wait for Clk_period;
		Addr <=  "00001111111011";
		Trees_din <= x"1401ce04";
		wait for Clk_period;
		Addr <=  "00001111111100";
		Trees_din <= x"fff71001";
		wait for Clk_period;
		Addr <=  "00001111111101";
		Trees_din <= x"0502dc04";
		wait for Clk_period;
		Addr <=  "00001111111110";
		Trees_din <= x"002c1001";
		wait for Clk_period;
		Addr <=  "00001111111111";
		Trees_din <= x"00041001";
		wait for Clk_period;
		Addr <=  "00010000000000";
		Trees_din <= x"01124608";
		wait for Clk_period;
		Addr <=  "00010000000001";
		Trees_din <= x"06ffd704";
		wait for Clk_period;
		Addr <=  "00010000000010";
		Trees_din <= x"0003101d";
		wait for Clk_period;
		Addr <=  "00010000000011";
		Trees_din <= x"ffd9101d";
		wait for Clk_period;
		Addr <=  "00010000000100";
		Trees_din <= x"040ebb04";
		wait for Clk_period;
		Addr <=  "00010000000101";
		Trees_din <= x"0028101d";
		wait for Clk_period;
		Addr <=  "00010000000110";
		Trees_din <= x"0006101d";
		wait for Clk_period;
		Addr <=  "00010000000111";
		Trees_din <= x"01037504";
		wait for Clk_period;
		Addr <=  "00010000001000";
		Trees_din <= x"ffe01039";
		wait for Clk_period;
		Addr <=  "00010000001001";
		Trees_din <= x"16007108";
		wait for Clk_period;
		Addr <=  "00010000001010";
		Trees_din <= x"15028704";
		wait for Clk_period;
		Addr <=  "00010000001011";
		Trees_din <= x"00131039";
		wait for Clk_period;
		Addr <=  "00010000001100";
		Trees_din <= x"ffe41039";
		wait for Clk_period;
		Addr <=  "00010000001101";
		Trees_din <= x"00211039";
		wait for Clk_period;
		Addr <=  "00010000001110";
		Trees_din <= x"01037504";
		wait for Clk_period;
		Addr <=  "00010000001111";
		Trees_din <= x"ffe21055";
		wait for Clk_period;
		Addr <=  "00010000010000";
		Trees_din <= x"07005404";
		wait for Clk_period;
		Addr <=  "00010000010001";
		Trees_din <= x"fff31055";
		wait for Clk_period;
		Addr <=  "00010000010010";
		Trees_din <= x"13023504";
		wait for Clk_period;
		Addr <=  "00010000010011";
		Trees_din <= x"00271055";
		wait for Clk_period;
		Addr <=  "00010000010100";
		Trees_din <= x"fffa1055";
		wait for Clk_period;
		Addr <=  "00010000010101";
		Trees_din <= x"01002704";
		wait for Clk_period;
		Addr <=  "00010000010110";
		Trees_din <= x"ffe01079";
		wait for Clk_period;
		Addr <=  "00010000010111";
		Trees_din <= x"07005404";
		wait for Clk_period;
		Addr <=  "00010000011000";
		Trees_din <= x"fff01079";
		wait for Clk_period;
		Addr <=  "00010000011001";
		Trees_din <= x"13023508";
		wait for Clk_period;
		Addr <=  "00010000011010";
		Trees_din <= x"1b010e04";
		wait for Clk_period;
		Addr <=  "00010000011011";
		Trees_din <= x"002f1079";
		wait for Clk_period;
		Addr <=  "00010000011100";
		Trees_din <= x"00091079";
		wait for Clk_period;
		Addr <=  "00010000011101";
		Trees_din <= x"fff91079";
		wait for Clk_period;
		Addr <=  "00010000011110";
		Trees_din <= x"01037504";
		wait for Clk_period;
		Addr <=  "00010000011111";
		Trees_din <= x"ffe61095";
		wait for Clk_period;
		Addr <=  "00010000100000";
		Trees_din <= x"0a015908";
		wait for Clk_period;
		Addr <=  "00010000100001";
		Trees_din <= x"0502dc04";
		wait for Clk_period;
		Addr <=  "00010000100010";
		Trees_din <= x"00291095";
		wait for Clk_period;
		Addr <=  "00010000100011";
		Trees_din <= x"fffe1095";
		wait for Clk_period;
		Addr <=  "00010000100100";
		Trees_din <= x"fff91095";
		wait for Clk_period;
		Addr <=  "00010000100101";
		Trees_din <= x"01037504";
		wait for Clk_period;
		Addr <=  "00010000100110";
		Trees_din <= x"ffe710b1";
		wait for Clk_period;
		Addr <=  "00010000100111";
		Trees_din <= x"16007108";
		wait for Clk_period;
		Addr <=  "00010000101000";
		Trees_din <= x"0b010504";
		wait for Clk_period;
		Addr <=  "00010000101001";
		Trees_din <= x"ffe910b1";
		wait for Clk_period;
		Addr <=  "00010000101010";
		Trees_din <= x"000f10b1";
		wait for Clk_period;
		Addr <=  "00010000101011";
		Trees_din <= x"001a10b1";
		wait for Clk_period;
		Addr <=  "00010000101100";
		Trees_din <= x"02029904";
		wait for Clk_period;
		Addr <=  "00010000101101";
		Trees_din <= x"ffeb10cd";
		wait for Clk_period;
		Addr <=  "00010000101110";
		Trees_din <= x"011cba08";
		wait for Clk_period;
		Addr <=  "00010000101111";
		Trees_din <= x"04067304";
		wait for Clk_period;
		Addr <=  "00010000110000";
		Trees_din <= x"000e10cd";
		wait for Clk_period;
		Addr <=  "00010000110001";
		Trees_din <= x"ffde10cd";
		wait for Clk_period;
		Addr <=  "00010000110010";
		Trees_din <= x"002610cd";
		wait for Clk_period;
		Addr <=  "00010000110011";
		Trees_din <= x"1103120c";
		wait for Clk_period;
		Addr <=  "00010000110100";
		Trees_din <= x"1101af08";
		wait for Clk_period;
		Addr <=  "00010000110101";
		Trees_din <= x"1402b504";
		wait for Clk_period;
		Addr <=  "00010000110110";
		Trees_din <= x"001910e9";
		wait for Clk_period;
		Addr <=  "00010000110111";
		Trees_din <= x"ffed10e9";
		wait for Clk_period;
		Addr <=  "00010000111000";
		Trees_din <= x"ffe110e9";
		wait for Clk_period;
		Addr <=  "00010000111001";
		Trees_din <= x"001610e9";
		wait for Clk_period;
		Addr <=  "00010000111010";
		Trees_din <= x"01037504";
		wait for Clk_period;
		Addr <=  "00010000111011";
		Trees_din <= x"ffe71105";
		wait for Clk_period;
		Addr <=  "00010000111100";
		Trees_din <= x"1c003004";
		wait for Clk_period;
		Addr <=  "00010000111101";
		Trees_din <= x"001c1105";
		wait for Clk_period;
		Addr <=  "00010000111110";
		Trees_din <= x"0a015904";
		wait for Clk_period;
		Addr <=  "00010000111111";
		Trees_din <= x"00101105";
		wait for Clk_period;
		Addr <=  "00010001000000";
		Trees_din <= x"ffee1105";
		wait for Clk_period;
		Addr <=  "00010001000001";
		Trees_din <= x"02097e08";
		wait for Clk_period;
		Addr <=  "00010001000010";
		Trees_din <= x"1b019a04";
		wait for Clk_period;
		Addr <=  "00010001000011";
		Trees_din <= x"ffdf1121";
		wait for Clk_period;
		Addr <=  "00010001000100";
		Trees_din <= x"00091121";
		wait for Clk_period;
		Addr <=  "00010001000101";
		Trees_din <= x"0b008804";
		wait for Clk_period;
		Addr <=  "00010001000110";
		Trees_din <= x"fff71121";
		wait for Clk_period;
		Addr <=  "00010001000111";
		Trees_din <= x"001e1121";
		wait for Clk_period;
		Addr <=  "00010001001000";
		Trees_din <= x"13fb9604";
		wait for Clk_period;
		Addr <=  "00010001001001";
		Trees_din <= x"ffee113d";
		wait for Clk_period;
		Addr <=  "00010001001010";
		Trees_din <= x"08005708";
		wait for Clk_period;
		Addr <=  "00010001001011";
		Trees_din <= x"1e006504";
		wait for Clk_period;
		Addr <=  "00010001001100";
		Trees_din <= x"fffe113d";
		wait for Clk_period;
		Addr <=  "00010001001101";
		Trees_din <= x"0024113d";
		wait for Clk_period;
		Addr <=  "00010001001110";
		Trees_din <= x"ffed113d";
		wait for Clk_period;
		Addr <=  "00010001001111";
		Trees_din <= x"01037504";
		wait for Clk_period;
		Addr <=  "00010001010000";
		Trees_din <= x"ffe71159";
		wait for Clk_period;
		Addr <=  "00010001010001";
		Trees_din <= x"1100e204";
		wait for Clk_period;
		Addr <=  "00010001010010";
		Trees_din <= x"fff71159";
		wait for Clk_period;
		Addr <=  "00010001010011";
		Trees_din <= x"011a8c04";
		wait for Clk_period;
		Addr <=  "00010001010100";
		Trees_din <= x"fffc1159";
		wait for Clk_period;
		Addr <=  "00010001010101";
		Trees_din <= x"00291159";
		wait for Clk_period;
		Addr <=  "00010001010110";
		Trees_din <= x"17004a0c";
		wait for Clk_period;
		Addr <=  "00010001010111";
		Trees_din <= x"011a8c08";
		wait for Clk_period;
		Addr <=  "00010001011000";
		Trees_din <= x"03fd1f04";
		wait for Clk_period;
		Addr <=  "00010001011001";
		Trees_din <= x"00081175";
		wait for Clk_period;
		Addr <=  "00010001011010";
		Trees_din <= x"ffe11175";
		wait for Clk_period;
		Addr <=  "00010001011011";
		Trees_din <= x"00301175";
		wait for Clk_period;
		Addr <=  "00010001011100";
		Trees_din <= x"ffed1175";
		wait for Clk_period;
		Addr <=  "00010001011101";
		Trees_din <= x"02097e08";
		wait for Clk_period;
		Addr <=  "00010001011110";
		Trees_din <= x"1b023d04";
		wait for Clk_period;
		Addr <=  "00010001011111";
		Trees_din <= x"ffe61191";
		wait for Clk_period;
		Addr <=  "00010001100000";
		Trees_din <= x"000a1191";
		wait for Clk_period;
		Addr <=  "00010001100001";
		Trees_din <= x"0b008804";
		wait for Clk_period;
		Addr <=  "00010001100010";
		Trees_din <= x"fff61191";
		wait for Clk_period;
		Addr <=  "00010001100011";
		Trees_din <= x"001c1191";
		wait for Clk_period;
		Addr <=  "00010001100100";
		Trees_din <= x"01037504";
		wait for Clk_period;
		Addr <=  "00010001100101";
		Trees_din <= x"ffe811ad";
		wait for Clk_period;
		Addr <=  "00010001100110";
		Trees_din <= x"1401ce04";
		wait for Clk_period;
		Addr <=  "00010001100111";
		Trees_din <= x"fff911ad";
		wait for Clk_period;
		Addr <=  "00010001101000";
		Trees_din <= x"1601fb04";
		wait for Clk_period;
		Addr <=  "00010001101001";
		Trees_din <= x"001e11ad";
		wait for Clk_period;
		Addr <=  "00010001101010";
		Trees_din <= x"000211ad";
		wait for Clk_period;
		Addr <=  "00010001101011";
		Trees_din <= x"02029904";
		wait for Clk_period;
		Addr <=  "00010001101100";
		Trees_din <= x"ffef11c9";
		wait for Clk_period;
		Addr <=  "00010001101101";
		Trees_din <= x"0efc6a04";
		wait for Clk_period;
		Addr <=  "00010001101110";
		Trees_din <= x"fff311c9";
		wait for Clk_period;
		Addr <=  "00010001101111";
		Trees_din <= x"07005704";
		wait for Clk_period;
		Addr <=  "00010001110000";
		Trees_din <= x"002011c9";
		wait for Clk_period;
		Addr <=  "00010001110001";
		Trees_din <= x"fffe11c9";
		wait for Clk_period;
		Addr <=  "00010001110010";
		Trees_din <= x"13fb9604";
		wait for Clk_period;
		Addr <=  "00010001110011";
		Trees_din <= x"fff011dd";
		wait for Clk_period;
		Addr <=  "00010001110100";
		Trees_din <= x"01081b04";
		wait for Clk_period;
		Addr <=  "00010001110101";
		Trees_din <= x"fff011dd";
		wait for Clk_period;
		Addr <=  "00010001110110";
		Trees_din <= x"001911dd";
		wait for Clk_period;
		Addr <=  "00010001110111";
		Trees_din <= x"17004a08";
		wait for Clk_period;
		Addr <=  "00010001111000";
		Trees_din <= x"010d0404";
		wait for Clk_period;
		Addr <=  "00010001111001";
		Trees_din <= x"ffeb11f1";
		wait for Clk_period;
		Addr <=  "00010001111010";
		Trees_din <= x"001f11f1";
		wait for Clk_period;
		Addr <=  "00010001111011";
		Trees_din <= x"ffef11f1";
		wait for Clk_period;
		Addr <=  "00010001111100";
		Trees_din <= x"19009508";
		wait for Clk_period;
		Addr <=  "00010001111101";
		Trees_din <= x"17004a04";
		wait for Clk_period;
		Addr <=  "00010001111110";
		Trees_din <= x"0020120d";
		wait for Clk_period;
		Addr <=  "00010001111111";
		Trees_din <= x"fff1120d";
		wait for Clk_period;
		Addr <=  "00010010000000";
		Trees_din <= x"16007104";
		wait for Clk_period;
		Addr <=  "00010010000001";
		Trees_din <= x"ffe7120d";
		wait for Clk_period;
		Addr <=  "00010010000010";
		Trees_din <= x"0007120d";
		wait for Clk_period;
		Addr <=  "00010010000011";
		Trees_din <= x"0bfda404";
		wait for Clk_period;
		Addr <=  "00010010000100";
		Trees_din <= x"00101221";
		wait for Clk_period;
		Addr <=  "00010010000101";
		Trees_din <= x"010d0404";
		wait for Clk_period;
		Addr <=  "00010010000110";
		Trees_din <= x"ffe21221";
		wait for Clk_period;
		Addr <=  "00010010000111";
		Trees_din <= x"000d1221";
		wait for Clk_period;
		Addr <=  "00010010001000";
		Trees_din <= x"02097e08";
		wait for Clk_period;
		Addr <=  "00010010001001";
		Trees_din <= x"1b019a04";
		wait for Clk_period;
		Addr <=  "00010010001010";
		Trees_din <= x"ffe6123d";
		wait for Clk_period;
		Addr <=  "00010010001011";
		Trees_din <= x"0007123d";
		wait for Clk_period;
		Addr <=  "00010010001100";
		Trees_din <= x"040ebb04";
		wait for Clk_period;
		Addr <=  "00010010001101";
		Trees_din <= x"0018123d";
		wait for Clk_period;
		Addr <=  "00010010001110";
		Trees_din <= x"fff7123d";
		wait for Clk_period;
		Addr <=  "00010010001111";
		Trees_din <= x"0bfda404";
		wait for Clk_period;
		Addr <=  "00010010010000";
		Trees_din <= x"000f1251";
		wait for Clk_period;
		Addr <=  "00010010010001";
		Trees_din <= x"010d0404";
		wait for Clk_period;
		Addr <=  "00010010010010";
		Trees_din <= x"ffe41251";
		wait for Clk_period;
		Addr <=  "00010010010011";
		Trees_din <= x"000c1251";
		wait for Clk_period;
		Addr <=  "00010010010100";
		Trees_din <= x"07005404";
		wait for Clk_period;
		Addr <=  "00010010010101";
		Trees_din <= x"fff11265";
		wait for Clk_period;
		Addr <=  "00010010010110";
		Trees_din <= x"08005704";
		wait for Clk_period;
		Addr <=  "00010010010111";
		Trees_din <= x"00161265";
		wait for Clk_period;
		Addr <=  "00010010011000";
		Trees_din <= x"fff01265";
		wait for Clk_period;
		Addr <=  "00010010011001";
		Trees_din <= x"1d00da08";
		wait for Clk_period;
		Addr <=  "00010010011010";
		Trees_din <= x"0f01cc04";
		wait for Clk_period;
		Addr <=  "00010010011011";
		Trees_din <= x"000b1279";
		wait for Clk_period;
		Addr <=  "00010010011100";
		Trees_din <= x"ffe61279";
		wait for Clk_period;
		Addr <=  "00010010011101";
		Trees_din <= x"000e1279";
		wait for Clk_period;
		Addr <=  "00010010011110";
		Trees_din <= x"1c003608";
		wait for Clk_period;
		Addr <=  "00010010011111";
		Trees_din <= x"16007104";
		wait for Clk_period;
		Addr <=  "00010010100000";
		Trees_din <= x"ffe91295";
		wait for Clk_period;
		Addr <=  "00010010100001";
		Trees_din <= x"00071295";
		wait for Clk_period;
		Addr <=  "00010010100010";
		Trees_din <= x"17004a04";
		wait for Clk_period;
		Addr <=  "00010010100011";
		Trees_din <= x"001d1295";
		wait for Clk_period;
		Addr <=  "00010010100100";
		Trees_din <= x"fff21295";
		wait for Clk_period;
		Addr <=  "00010010100101";
		Trees_din <= x"1d00da08";
		wait for Clk_period;
		Addr <=  "00010010100110";
		Trees_din <= x"05027104";
		wait for Clk_period;
		Addr <=  "00010010100111";
		Trees_din <= x"000a12a9";
		wait for Clk_period;
		Addr <=  "00010010101000";
		Trees_din <= x"ffe712a9";
		wait for Clk_period;
		Addr <=  "00010010101001";
		Trees_din <= x"000e12a9";
		wait for Clk_period;
		Addr <=  "00010010101010";
		Trees_din <= x"02097e08";
		wait for Clk_period;
		Addr <=  "00010010101011";
		Trees_din <= x"19009504";
		wait for Clk_period;
		Addr <=  "00010010101100";
		Trees_din <= x"000612c5";
		wait for Clk_period;
		Addr <=  "00010010101101";
		Trees_din <= x"ffe812c5";
		wait for Clk_period;
		Addr <=  "00010010101110";
		Trees_din <= x"1300c004";
		wait for Clk_period;
		Addr <=  "00010010101111";
		Trees_din <= x"001412c5";
		wait for Clk_period;
		Addr <=  "00010010110000";
		Trees_din <= x"fffb12c5";
		wait for Clk_period;
		Addr <=  "00010010110001";
		Trees_din <= x"1d00da08";
		wait for Clk_period;
		Addr <=  "00010010110010";
		Trees_din <= x"0f01cc04";
		wait for Clk_period;
		Addr <=  "00010010110011";
		Trees_din <= x"000a12d9";
		wait for Clk_period;
		Addr <=  "00010010110100";
		Trees_din <= x"ffe812d9";
		wait for Clk_period;
		Addr <=  "00010010110101";
		Trees_din <= x"000d12d9";
		wait for Clk_period;
		Addr <=  "00010010110110";
		Trees_din <= x"10021408";
		wait for Clk_period;
		Addr <=  "00010010110111";
		Trees_din <= x"0f013304";
		wait for Clk_period;
		Addr <=  "00010010111000";
		Trees_din <= x"000612ed";
		wait for Clk_period;
		Addr <=  "00010010111001";
		Trees_din <= x"ffe712ed";
		wait for Clk_period;
		Addr <=  "00010010111010";
		Trees_din <= x"000c12ed";
		wait for Clk_period;
		Addr <=  "00010010111011";
		Trees_din <= x"02097e08";
		wait for Clk_period;
		Addr <=  "00010010111100";
		Trees_din <= x"1b019a04";
		wait for Clk_period;
		Addr <=  "00010010111101";
		Trees_din <= x"ffe91309";
		wait for Clk_period;
		Addr <=  "00010010111110";
		Trees_din <= x"00061309";
		wait for Clk_period;
		Addr <=  "00010010111111";
		Trees_din <= x"1300c004";
		wait for Clk_period;
		Addr <=  "00010011000000";
		Trees_din <= x"00141309";
		wait for Clk_period;
		Addr <=  "00010011000001";
		Trees_din <= x"fffb1309";
		wait for Clk_period;
		Addr <=  "00010011000010";
		Trees_din <= x"0bfda404";
		wait for Clk_period;
		Addr <=  "00010011000011";
		Trees_din <= x"000d1325";
		wait for Clk_period;
		Addr <=  "00010011000100";
		Trees_din <= x"15044908";
		wait for Clk_period;
		Addr <=  "00010011000101";
		Trees_din <= x"02097e04";
		wait for Clk_period;
		Addr <=  "00010011000110";
		Trees_din <= x"fff41325";
		wait for Clk_period;
		Addr <=  "00010011000111";
		Trees_din <= x"00171325";
		wait for Clk_period;
		Addr <=  "00010011001000";
		Trees_din <= x"ffe51325";
		wait for Clk_period;
		Addr <=  "00010011001001";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  4
        -----------
		Addr <=  "00000000000000";
		Trees_din <= x"020d6230";
		wait for Clk_period;
		Addr <=  "00000000000001";
		Trees_din <= x"0209d118";
		wait for Clk_period;
		Addr <=  "00000000000010";
		Trees_din <= x"02072404";
		wait for Clk_period;
		Addr <=  "00000000000011";
		Trees_din <= x"ff4e008d";
		wait for Clk_period;
		Addr <=  "00000000000100";
		Trees_din <= x"00019008";
		wait for Clk_period;
		Addr <=  "00000000000101";
		Trees_din <= x"1603f604";
		wait for Clk_period;
		Addr <=  "00000000000110";
		Trees_din <= x"ff51008d";
		wait for Clk_period;
		Addr <=  "00000000000111";
		Trees_din <= x"0027008d";
		wait for Clk_period;
		Addr <=  "00000000001000";
		Trees_din <= x"000c1008";
		wait for Clk_period;
		Addr <=  "00000000001001";
		Trees_din <= x"0506ce04";
		wait for Clk_period;
		Addr <=  "00000000001010";
		Trees_din <= x"0275008d";
		wait for Clk_period;
		Addr <=  "00000000001011";
		Trees_din <= x"ffe5008d";
		wait for Clk_period;
		Addr <=  "00000000001100";
		Trees_din <= x"ff61008d";
		wait for Clk_period;
		Addr <=  "00000000001101";
		Trees_din <= x"00f0ae08";
		wait for Clk_period;
		Addr <=  "00000000001110";
		Trees_din <= x"10fd9004";
		wait for Clk_period;
		Addr <=  "00000000001111";
		Trees_din <= x"0000008d";
		wait for Clk_period;
		Addr <=  "00000000010000";
		Trees_din <= x"ff53008d";
		wait for Clk_period;
		Addr <=  "00000000010001";
		Trees_din <= x"000c100c";
		wait for Clk_period;
		Addr <=  "00000000010010";
		Trees_din <= x"06fc4208";
		wait for Clk_period;
		Addr <=  "00000000010011";
		Trees_din <= x"00026604";
		wait for Clk_period;
		Addr <=  "00000000010100";
		Trees_din <= x"ff89008d";
		wait for Clk_period;
		Addr <=  "00000000010101";
		Trees_din <= x"013c008d";
		wait for Clk_period;
		Addr <=  "00000000010110";
		Trees_din <= x"038d008d";
		wait for Clk_period;
		Addr <=  "00000000010111";
		Trees_din <= x"ff85008d";
		wait for Clk_period;
		Addr <=  "00000000011000";
		Trees_din <= x"011a8c10";
		wait for Clk_period;
		Addr <=  "00000000011001";
		Trees_din <= x"06175708";
		wait for Clk_period;
		Addr <=  "00000000011010";
		Trees_din <= x"05150f04";
		wait for Clk_period;
		Addr <=  "00000000011011";
		Trees_din <= x"041f008d";
		wait for Clk_period;
		Addr <=  "00000000011100";
		Trees_din <= x"ff75008d";
		wait for Clk_period;
		Addr <=  "00000000011101";
		Trees_din <= x"061cb504";
		wait for Clk_period;
		Addr <=  "00000000011110";
		Trees_din <= x"0027008d";
		wait for Clk_period;
		Addr <=  "00000000011111";
		Trees_din <= x"ff6e008d";
		wait for Clk_period;
		Addr <=  "00000000100000";
		Trees_din <= x"021ddb04";
		wait for Clk_period;
		Addr <=  "00000000100001";
		Trees_din <= x"ff56008d";
		wait for Clk_period;
		Addr <=  "00000000100010";
		Trees_din <= x"0280008d";
		wait for Clk_period;
		Addr <=  "00000000100011";
		Trees_din <= x"020b1e2c";
		wait for Clk_period;
		Addr <=  "00000000100100";
		Trees_din <= x"02072414";
		wait for Clk_period;
		Addr <=  "00000000100101";
		Trees_din <= x"1b03ff0c";
		wait for Clk_period;
		Addr <=  "00000000100110";
		Trees_din <= x"14040004";
		wait for Clk_period;
		Addr <=  "00000000100111";
		Trees_din <= x"ff550131";
		wait for Clk_period;
		Addr <=  "00000000101000";
		Trees_din <= x"02030104";
		wait for Clk_period;
		Addr <=  "00000000101001";
		Trees_din <= x"ff5f0131";
		wait for Clk_period;
		Addr <=  "00000000101010";
		Trees_din <= x"00800131";
		wait for Clk_period;
		Addr <=  "00000000101011";
		Trees_din <= x"0a000104";
		wait for Clk_period;
		Addr <=  "00000000101100";
		Trees_din <= x"00340131";
		wait for Clk_period;
		Addr <=  "00000000101101";
		Trees_din <= x"ff780131";
		wait for Clk_period;
		Addr <=  "00000000101110";
		Trees_din <= x"00fc1104";
		wait for Clk_period;
		Addr <=  "00000000101111";
		Trees_din <= x"ff570131";
		wait for Clk_period;
		Addr <=  "00000000110000";
		Trees_din <= x"000c1010";
		wait for Clk_period;
		Addr <=  "00000000110001";
		Trees_din <= x"05054b08";
		wait for Clk_period;
		Addr <=  "00000000110010";
		Trees_din <= x"04009e04";
		wait for Clk_period;
		Addr <=  "00000000110011";
		Trees_din <= x"01f20131";
		wait for Clk_period;
		Addr <=  "00000000110100";
		Trees_din <= x"ff840131";
		wait for Clk_period;
		Addr <=  "00000000110101";
		Trees_din <= x"10028704";
		wait for Clk_period;
		Addr <=  "00000000110110";
		Trees_din <= x"ff6b0131";
		wait for Clk_period;
		Addr <=  "00000000110111";
		Trees_din <= x"00a90131";
		wait for Clk_period;
		Addr <=  "00000000111000";
		Trees_din <= x"ff690131";
		wait for Clk_period;
		Addr <=  "00000000111001";
		Trees_din <= x"0116f11c";
		wait for Clk_period;
		Addr <=  "00000000111010";
		Trees_din <= x"06175714";
		wait for Clk_period;
		Addr <=  "00000000111011";
		Trees_din <= x"05119e0c";
		wait for Clk_period;
		Addr <=  "00000000111100";
		Trees_din <= x"000c1008";
		wait for Clk_period;
		Addr <=  "00000000111101";
		Trees_din <= x"050e0404";
		wait for Clk_period;
		Addr <=  "00000000111110";
		Trees_din <= x"01a80131";
		wait for Clk_period;
		Addr <=  "00000000111111";
		Trees_din <= x"00ae0131";
		wait for Clk_period;
		Addr <=  "00000001000000";
		Trees_din <= x"ff940131";
		wait for Clk_period;
		Addr <=  "00000001000001";
		Trees_din <= x"08005904";
		wait for Clk_period;
		Addr <=  "00000001000010";
		Trees_din <= x"ff6e0131";
		wait for Clk_period;
		Addr <=  "00000001000011";
		Trees_din <= x"00340131";
		wait for Clk_period;
		Addr <=  "00000001000100";
		Trees_din <= x"1b035a04";
		wait for Clk_period;
		Addr <=  "00000001000101";
		Trees_din <= x"ff6c0131";
		wait for Clk_period;
		Addr <=  "00000001000110";
		Trees_din <= x"003c0131";
		wait for Clk_period;
		Addr <=  "00000001000111";
		Trees_din <= x"021b0604";
		wait for Clk_period;
		Addr <=  "00000001001000";
		Trees_din <= x"ff580131";
		wait for Clk_period;
		Addr <=  "00000001001001";
		Trees_din <= x"0ffeb904";
		wait for Clk_period;
		Addr <=  "00000001001010";
		Trees_din <= x"00230131";
		wait for Clk_period;
		Addr <=  "00000001001011";
		Trees_din <= x"01a80131";
		wait for Clk_period;
		Addr <=  "00000001001100";
		Trees_din <= x"020b1e2c";
		wait for Clk_period;
		Addr <=  "00000001001101";
		Trees_din <= x"02072418";
		wait for Clk_period;
		Addr <=  "00000001001110";
		Trees_din <= x"02030104";
		wait for Clk_period;
		Addr <=  "00000001001111";
		Trees_din <= x"ff5901cd";
		wait for Clk_period;
		Addr <=  "00000001010000";
		Trees_din <= x"1603fa10";
		wait for Clk_period;
		Addr <=  "00000001010001";
		Trees_din <= x"0a000108";
		wait for Clk_period;
		Addr <=  "00000001010010";
		Trees_din <= x"0d018a04";
		wait for Clk_period;
		Addr <=  "00000001010011";
		Trees_din <= x"ff6d01cd";
		wait for Clk_period;
		Addr <=  "00000001010100";
		Trees_din <= x"00a201cd";
		wait for Clk_period;
		Addr <=  "00000001010101";
		Trees_din <= x"02031d04";
		wait for Clk_period;
		Addr <=  "00000001010110";
		Trees_din <= x"ffb001cd";
		wait for Clk_period;
		Addr <=  "00000001010111";
		Trees_din <= x"ff5d01cd";
		wait for Clk_period;
		Addr <=  "00000001011000";
		Trees_din <= x"007f01cd";
		wait for Clk_period;
		Addr <=  "00000001011001";
		Trees_din <= x"00fc1104";
		wait for Clk_period;
		Addr <=  "00000001011010";
		Trees_din <= x"ff5c01cd";
		wait for Clk_period;
		Addr <=  "00000001011011";
		Trees_din <= x"000c100c";
		wait for Clk_period;
		Addr <=  "00000001011100";
		Trees_din <= x"05098d08";
		wait for Clk_period;
		Addr <=  "00000001011101";
		Trees_din <= x"04009e04";
		wait for Clk_period;
		Addr <=  "00000001011110";
		Trees_din <= x"012f01cd";
		wait for Clk_period;
		Addr <=  "00000001011111";
		Trees_din <= x"ff8701cd";
		wait for Clk_period;
		Addr <=  "00000001100000";
		Trees_din <= x"ff7d01cd";
		wait for Clk_period;
		Addr <=  "00000001100001";
		Trees_din <= x"ff7101cd";
		wait for Clk_period;
		Addr <=  "00000001100010";
		Trees_din <= x"011cba1c";
		wait for Clk_period;
		Addr <=  "00000001100011";
		Trees_din <= x"06175714";
		wait for Clk_period;
		Addr <=  "00000001100100";
		Trees_din <= x"05119e0c";
		wait for Clk_period;
		Addr <=  "00000001100101";
		Trees_din <= x"020f1908";
		wait for Clk_period;
		Addr <=  "00000001100110";
		Trees_din <= x"00f0ae04";
		wait for Clk_period;
		Addr <=  "00000001100111";
		Trees_din <= x"ff7c01cd";
		wait for Clk_period;
		Addr <=  "00000001101000";
		Trees_din <= x"011501cd";
		wait for Clk_period;
		Addr <=  "00000001101001";
		Trees_din <= x"013401cd";
		wait for Clk_period;
		Addr <=  "00000001101010";
		Trees_din <= x"040db704";
		wait for Clk_period;
		Addr <=  "00000001101011";
		Trees_din <= x"ff7301cd";
		wait for Clk_period;
		Addr <=  "00000001101100";
		Trees_din <= x"00b701cd";
		wait for Clk_period;
		Addr <=  "00000001101101";
		Trees_din <= x"0a000f04";
		wait for Clk_period;
		Addr <=  "00000001101110";
		Trees_din <= x"003001cd";
		wait for Clk_period;
		Addr <=  "00000001101111";
		Trees_din <= x"ff6f01cd";
		wait for Clk_period;
		Addr <=  "00000001110000";
		Trees_din <= x"050e0404";
		wait for Clk_period;
		Addr <=  "00000001110001";
		Trees_din <= x"ff6301cd";
		wait for Clk_period;
		Addr <=  "00000001110010";
		Trees_din <= x"003e01cd";
		wait for Clk_period;
		Addr <=  "00000001110011";
		Trees_din <= x"020b1e30";
		wait for Clk_period;
		Addr <=  "00000001110100";
		Trees_din <= x"02072418";
		wait for Clk_period;
		Addr <=  "00000001110101";
		Trees_din <= x"02030104";
		wait for Clk_period;
		Addr <=  "00000001110110";
		Trees_din <= x"ff5c0271";
		wait for Clk_period;
		Addr <=  "00000001110111";
		Trees_din <= x"1603fa10";
		wait for Clk_period;
		Addr <=  "00000001111000";
		Trees_din <= x"0a000108";
		wait for Clk_period;
		Addr <=  "00000001111001";
		Trees_din <= x"0d018a04";
		wait for Clk_period;
		Addr <=  "00000001111010";
		Trees_din <= x"ff740271";
		wait for Clk_period;
		Addr <=  "00000001111011";
		Trees_din <= x"00900271";
		wait for Clk_period;
		Addr <=  "00000001111100";
		Trees_din <= x"02031d04";
		wait for Clk_period;
		Addr <=  "00000001111101";
		Trees_din <= x"ffbe0271";
		wait for Clk_period;
		Addr <=  "00000001111110";
		Trees_din <= x"ff620271";
		wait for Clk_period;
		Addr <=  "00000001111111";
		Trees_din <= x"00710271";
		wait for Clk_period;
		Addr <=  "00000010000000";
		Trees_din <= x"00fc1104";
		wait for Clk_period;
		Addr <=  "00000010000001";
		Trees_din <= x"ff610271";
		wait for Clk_period;
		Addr <=  "00000010000010";
		Trees_din <= x"000c1010";
		wait for Clk_period;
		Addr <=  "00000010000011";
		Trees_din <= x"05054b08";
		wait for Clk_period;
		Addr <=  "00000010000100";
		Trees_din <= x"04009e04";
		wait for Clk_period;
		Addr <=  "00000010000101";
		Trees_din <= x"010d0271";
		wait for Clk_period;
		Addr <=  "00000010000110";
		Trees_din <= x"ff910271";
		wait for Clk_period;
		Addr <=  "00000010000111";
		Trees_din <= x"10028704";
		wait for Clk_period;
		Addr <=  "00000010001000";
		Trees_din <= x"ff6d0271";
		wait for Clk_period;
		Addr <=  "00000010001001";
		Trees_din <= x"00820271";
		wait for Clk_period;
		Addr <=  "00000010001010";
		Trees_din <= x"ff780271";
		wait for Clk_period;
		Addr <=  "00000010001011";
		Trees_din <= x"011cba1c";
		wait for Clk_period;
		Addr <=  "00000010001100";
		Trees_din <= x"06175714";
		wait for Clk_period;
		Addr <=  "00000010001101";
		Trees_din <= x"05119e0c";
		wait for Clk_period;
		Addr <=  "00000010001110";
		Trees_din <= x"000c1008";
		wait for Clk_period;
		Addr <=  "00000010001111";
		Trees_din <= x"0113b304";
		wait for Clk_period;
		Addr <=  "00000010010000";
		Trees_din <= x"00f60271";
		wait for Clk_period;
		Addr <=  "00000010010001";
		Trees_din <= x"00830271";
		wait for Clk_period;
		Addr <=  "00000010010010";
		Trees_din <= x"ff970271";
		wait for Clk_period;
		Addr <=  "00000010010011";
		Trees_din <= x"030a2c04";
		wait for Clk_period;
		Addr <=  "00000010010100";
		Trees_din <= x"ff7a0271";
		wait for Clk_period;
		Addr <=  "00000010010101";
		Trees_din <= x"009c0271";
		wait for Clk_period;
		Addr <=  "00000010010110";
		Trees_din <= x"1b035a04";
		wait for Clk_period;
		Addr <=  "00000010010111";
		Trees_din <= x"ff760271";
		wait for Clk_period;
		Addr <=  "00000010011000";
		Trees_din <= x"00330271";
		wait for Clk_period;
		Addr <=  "00000010011001";
		Trees_din <= x"050e0404";
		wait for Clk_period;
		Addr <=  "00000010011010";
		Trees_din <= x"ff690271";
		wait for Clk_period;
		Addr <=  "00000010011011";
		Trees_din <= x"00330271";
		wait for Clk_period;
		Addr <=  "00000010011100";
		Trees_din <= x"020b1e30";
		wait for Clk_period;
		Addr <=  "00000010011101";
		Trees_din <= x"02072418";
		wait for Clk_period;
		Addr <=  "00000010011110";
		Trees_din <= x"02030104";
		wait for Clk_period;
		Addr <=  "00000010011111";
		Trees_din <= x"ff5f0315";
		wait for Clk_period;
		Addr <=  "00000010100000";
		Trees_din <= x"14040010";
		wait for Clk_period;
		Addr <=  "00000010100001";
		Trees_din <= x"0a000108";
		wait for Clk_period;
		Addr <=  "00000010100010";
		Trees_din <= x"13028704";
		wait for Clk_period;
		Addr <=  "00000010100011";
		Trees_din <= x"ff790315";
		wait for Clk_period;
		Addr <=  "00000010100100";
		Trees_din <= x"00800315";
		wait for Clk_period;
		Addr <=  "00000010100101";
		Trees_din <= x"0bf98004";
		wait for Clk_period;
		Addr <=  "00000010100110";
		Trees_din <= x"ffd20315";
		wait for Clk_period;
		Addr <=  "00000010100111";
		Trees_din <= x"ff660315";
		wait for Clk_period;
		Addr <=  "00000010101000";
		Trees_din <= x"00680315";
		wait for Clk_period;
		Addr <=  "00000010101001";
		Trees_din <= x"00fc1104";
		wait for Clk_period;
		Addr <=  "00000010101010";
		Trees_din <= x"ff650315";
		wait for Clk_period;
		Addr <=  "00000010101011";
		Trees_din <= x"000c1010";
		wait for Clk_period;
		Addr <=  "00000010101100";
		Trees_din <= x"05054b08";
		wait for Clk_period;
		Addr <=  "00000010101101";
		Trees_din <= x"04009e04";
		wait for Clk_period;
		Addr <=  "00000010101110";
		Trees_din <= x"00e10315";
		wait for Clk_period;
		Addr <=  "00000010101111";
		Trees_din <= x"ff960315";
		wait for Clk_period;
		Addr <=  "00000010110000";
		Trees_din <= x"10028704";
		wait for Clk_period;
		Addr <=  "00000010110001";
		Trees_din <= x"ff720315";
		wait for Clk_period;
		Addr <=  "00000010110010";
		Trees_din <= x"006f0315";
		wait for Clk_period;
		Addr <=  "00000010110011";
		Trees_din <= x"ff800315";
		wait for Clk_period;
		Addr <=  "00000010110100";
		Trees_din <= x"011fa020";
		wait for Clk_period;
		Addr <=  "00000010110101";
		Trees_din <= x"020f1914";
		wait for Clk_period;
		Addr <=  "00000010110110";
		Trees_din <= x"00f0ae08";
		wait for Clk_period;
		Addr <=  "00000010110111";
		Trees_din <= x"0d03db04";
		wait for Clk_period;
		Addr <=  "00000010111000";
		Trees_din <= x"ff5f0315";
		wait for Clk_period;
		Addr <=  "00000010111001";
		Trees_din <= x"00290315";
		wait for Clk_period;
		Addr <=  "00000010111010";
		Trees_din <= x"04081e08";
		wait for Clk_period;
		Addr <=  "00000010111011";
		Trees_din <= x"000c1004";
		wait for Clk_period;
		Addr <=  "00000010111100";
		Trees_din <= x"00ce0315";
		wait for Clk_period;
		Addr <=  "00000010111101";
		Trees_din <= x"ffa10315";
		wait for Clk_period;
		Addr <=  "00000010111110";
		Trees_din <= x"ff780315";
		wait for Clk_period;
		Addr <=  "00000010111111";
		Trees_din <= x"061cb508";
		wait for Clk_period;
		Addr <=  "00000011000000";
		Trees_din <= x"0515e904";
		wait for Clk_period;
		Addr <=  "00000011000001";
		Trees_din <= x"00da0315";
		wait for Clk_period;
		Addr <=  "00000011000010";
		Trees_din <= x"fff60315";
		wait for Clk_period;
		Addr <=  "00000011000011";
		Trees_din <= x"ff950315";
		wait for Clk_period;
		Addr <=  "00000011000100";
		Trees_din <= x"ff6e0315";
		wait for Clk_period;
		Addr <=  "00000011000101";
		Trees_din <= x"020b1e24";
		wait for Clk_period;
		Addr <=  "00000011000110";
		Trees_din <= x"02056d0c";
		wait for Clk_period;
		Addr <=  "00000011000111";
		Trees_din <= x"14040004";
		wait for Clk_period;
		Addr <=  "00000011001000";
		Trees_din <= x"ff6203b1";
		wait for Clk_period;
		Addr <=  "00000011001001";
		Trees_din <= x"03fbeb04";
		wait for Clk_period;
		Addr <=  "00000011001010";
		Trees_din <= x"006703b1";
		wait for Clk_period;
		Addr <=  "00000011001011";
		Trees_din <= x"ff7703b1";
		wait for Clk_period;
		Addr <=  "00000011001100";
		Trees_din <= x"00fa7604";
		wait for Clk_period;
		Addr <=  "00000011001101";
		Trees_din <= x"ff6603b1";
		wait for Clk_period;
		Addr <=  "00000011001110";
		Trees_din <= x"000cbc10";
		wait for Clk_period;
		Addr <=  "00000011001111";
		Trees_din <= x"05054b08";
		wait for Clk_period;
		Addr <=  "00000011010000";
		Trees_din <= x"04009e04";
		wait for Clk_period;
		Addr <=  "00000011010001";
		Trees_din <= x"00ce03b1";
		wait for Clk_period;
		Addr <=  "00000011010010";
		Trees_din <= x"ff9303b1";
		wait for Clk_period;
		Addr <=  "00000011010011";
		Trees_din <= x"08004e04";
		wait for Clk_period;
		Addr <=  "00000011010100";
		Trees_din <= x"003b03b1";
		wait for Clk_period;
		Addr <=  "00000011010101";
		Trees_din <= x"ff6e03b1";
		wait for Clk_period;
		Addr <=  "00000011010110";
		Trees_din <= x"ff7603b1";
		wait for Clk_period;
		Addr <=  "00000011010111";
		Trees_din <= x"0116f120";
		wait for Clk_period;
		Addr <=  "00000011011000";
		Trees_din <= x"020f1914";
		wait for Clk_period;
		Addr <=  "00000011011001";
		Trees_din <= x"00f0ae08";
		wait for Clk_period;
		Addr <=  "00000011011010";
		Trees_din <= x"0d03b004";
		wait for Clk_period;
		Addr <=  "00000011011011";
		Trees_din <= x"ff6a03b1";
		wait for Clk_period;
		Addr <=  "00000011011100";
		Trees_din <= x"001703b1";
		wait for Clk_period;
		Addr <=  "00000011011101";
		Trees_din <= x"04081e08";
		wait for Clk_period;
		Addr <=  "00000011011110";
		Trees_din <= x"0d03e704";
		wait for Clk_period;
		Addr <=  "00000011011111";
		Trees_din <= x"00bc03b1";
		wait for Clk_period;
		Addr <=  "00000011100000";
		Trees_din <= x"ffd503b1";
		wait for Clk_period;
		Addr <=  "00000011100001";
		Trees_din <= x"ff8603b1";
		wait for Clk_period;
		Addr <=  "00000011100010";
		Trees_din <= x"061cb508";
		wait for Clk_period;
		Addr <=  "00000011100011";
		Trees_din <= x"05150f04";
		wait for Clk_period;
		Addr <=  "00000011100100";
		Trees_din <= x"00c703b1";
		wait for Clk_period;
		Addr <=  "00000011100101";
		Trees_din <= x"ffab03b1";
		wait for Clk_period;
		Addr <=  "00000011100110";
		Trees_din <= x"ffab03b1";
		wait for Clk_period;
		Addr <=  "00000011100111";
		Trees_din <= x"021b0604";
		wait for Clk_period;
		Addr <=  "00000011101000";
		Trees_din <= x"ff6803b1";
		wait for Clk_period;
		Addr <=  "00000011101001";
		Trees_din <= x"0ffeb904";
		wait for Clk_period;
		Addr <=  "00000011101010";
		Trees_din <= x"000103b1";
		wait for Clk_period;
		Addr <=  "00000011101011";
		Trees_din <= x"00c703b1";
		wait for Clk_period;
		Addr <=  "00000011101100";
		Trees_din <= x"020b1e24";
		wait for Clk_period;
		Addr <=  "00000011101101";
		Trees_din <= x"02056d0c";
		wait for Clk_period;
		Addr <=  "00000011101110";
		Trees_din <= x"14040004";
		wait for Clk_period;
		Addr <=  "00000011101111";
		Trees_din <= x"ff640455";
		wait for Clk_period;
		Addr <=  "00000011110000";
		Trees_din <= x"02030104";
		wait for Clk_period;
		Addr <=  "00000011110001";
		Trees_din <= x"ff7e0455";
		wait for Clk_period;
		Addr <=  "00000011110010";
		Trees_din <= x"006a0455";
		wait for Clk_period;
		Addr <=  "00000011110011";
		Trees_din <= x"00fa7604";
		wait for Clk_period;
		Addr <=  "00000011110100";
		Trees_din <= x"ff6a0455";
		wait for Clk_period;
		Addr <=  "00000011110101";
		Trees_din <= x"000cbc10";
		wait for Clk_period;
		Addr <=  "00000011110110";
		Trees_din <= x"05054b08";
		wait for Clk_period;
		Addr <=  "00000011110111";
		Trees_din <= x"04009e04";
		wait for Clk_period;
		Addr <=  "00000011111000";
		Trees_din <= x"00b50455";
		wait for Clk_period;
		Addr <=  "00000011111001";
		Trees_din <= x"ff970455";
		wait for Clk_period;
		Addr <=  "00000011111010";
		Trees_din <= x"08004e04";
		wait for Clk_period;
		Addr <=  "00000011111011";
		Trees_din <= x"00380455";
		wait for Clk_period;
		Addr <=  "00000011111100";
		Trees_din <= x"ff740455";
		wait for Clk_period;
		Addr <=  "00000011111101";
		Trees_din <= x"ff7d0455";
		wait for Clk_period;
		Addr <=  "00000011111110";
		Trees_din <= x"0113b320";
		wait for Clk_period;
		Addr <=  "00000011111111";
		Trees_din <= x"050e0414";
		wait for Clk_period;
		Addr <=  "00000100000000";
		Trees_din <= x"0617570c";
		wait for Clk_period;
		Addr <=  "00000100000001";
		Trees_din <= x"020f1908";
		wait for Clk_period;
		Addr <=  "00000100000010";
		Trees_din <= x"04081e04";
		wait for Clk_period;
		Addr <=  "00000100000011";
		Trees_din <= x"00910455";
		wait for Clk_period;
		Addr <=  "00000100000100";
		Trees_din <= x"ff860455";
		wait for Clk_period;
		Addr <=  "00000100000101";
		Trees_din <= x"00ba0455";
		wait for Clk_period;
		Addr <=  "00000100000110";
		Trees_din <= x"0d034004";
		wait for Clk_period;
		Addr <=  "00000100000111";
		Trees_din <= x"ffa20455";
		wait for Clk_period;
		Addr <=  "00000100001000";
		Trees_din <= x"00300455";
		wait for Clk_period;
		Addr <=  "00000100001001";
		Trees_din <= x"02117804";
		wait for Clk_period;
		Addr <=  "00000100001010";
		Trees_din <= x"ff820455";
		wait for Clk_period;
		Addr <=  "00000100001011";
		Trees_din <= x"0a00b304";
		wait for Clk_period;
		Addr <=  "00000100001100";
		Trees_din <= x"00730455";
		wait for Clk_period;
		Addr <=  "00000100001101";
		Trees_din <= x"001f0455";
		wait for Clk_period;
		Addr <=  "00000100001110";
		Trees_din <= x"021b0608";
		wait for Clk_period;
		Addr <=  "00000100001111";
		Trees_din <= x"02160e04";
		wait for Clk_period;
		Addr <=  "00000100010000";
		Trees_din <= x"ff660455";
		wait for Clk_period;
		Addr <=  "00000100010001";
		Trees_din <= x"fff10455";
		wait for Clk_period;
		Addr <=  "00000100010010";
		Trees_din <= x"0ffeb904";
		wait for Clk_period;
		Addr <=  "00000100010011";
		Trees_din <= x"fffd0455";
		wait for Clk_period;
		Addr <=  "00000100010100";
		Trees_din <= x"00b80455";
		wait for Clk_period;
		Addr <=  "00000100010101";
		Trees_din <= x"020b1e2c";
		wait for Clk_period;
		Addr <=  "00000100010110";
		Trees_din <= x"02056d0c";
		wait for Clk_period;
		Addr <=  "00000100010111";
		Trees_din <= x"14040004";
		wait for Clk_period;
		Addr <=  "00000100011000";
		Trees_din <= x"ff6604f9";
		wait for Clk_period;
		Addr <=  "00000100011001";
		Trees_din <= x"0a000704";
		wait for Clk_period;
		Addr <=  "00000100011010";
		Trees_din <= x"ff8304f9";
		wait for Clk_period;
		Addr <=  "00000100011011";
		Trees_din <= x"006a04f9";
		wait for Clk_period;
		Addr <=  "00000100011100";
		Trees_din <= x"00fa7604";
		wait for Clk_period;
		Addr <=  "00000100011101";
		Trees_din <= x"ff6d04f9";
		wait for Clk_period;
		Addr <=  "00000100011110";
		Trees_din <= x"06fe6f0c";
		wait for Clk_period;
		Addr <=  "00000100011111";
		Trees_din <= x"0a000004";
		wait for Clk_period;
		Addr <=  "00000100100000";
		Trees_din <= x"009904f9";
		wait for Clk_period;
		Addr <=  "00000100100001";
		Trees_din <= x"02083604";
		wait for Clk_period;
		Addr <=  "00000100100010";
		Trees_din <= x"ff7204f9";
		wait for Clk_period;
		Addr <=  "00000100100011";
		Trees_din <= x"001804f9";
		wait for Clk_period;
		Addr <=  "00000100100100";
		Trees_din <= x"08005708";
		wait for Clk_period;
		Addr <=  "00000100100101";
		Trees_din <= x"0a008c04";
		wait for Clk_period;
		Addr <=  "00000100100110";
		Trees_din <= x"005004f9";
		wait for Clk_period;
		Addr <=  "00000100100111";
		Trees_din <= x"ffc104f9";
		wait for Clk_period;
		Addr <=  "00000100101000";
		Trees_din <= x"1b01d304";
		wait for Clk_period;
		Addr <=  "00000100101001";
		Trees_din <= x"002804f9";
		wait for Clk_period;
		Addr <=  "00000100101010";
		Trees_din <= x"010f04f9";
		wait for Clk_period;
		Addr <=  "00000100101011";
		Trees_din <= x"011fa024";
		wait for Clk_period;
		Addr <=  "00000100101100";
		Trees_din <= x"020f1914";
		wait for Clk_period;
		Addr <=  "00000100101101";
		Trees_din <= x"00f0ae08";
		wait for Clk_period;
		Addr <=  "00000100101110";
		Trees_din <= x"08005904";
		wait for Clk_period;
		Addr <=  "00000100101111";
		Trees_din <= x"ff7004f9";
		wait for Clk_period;
		Addr <=  "00000100110000";
		Trees_din <= x"001f04f9";
		wait for Clk_period;
		Addr <=  "00000100110001";
		Trees_din <= x"06f98e04";
		wait for Clk_period;
		Addr <=  "00000100110010";
		Trees_din <= x"ff8d04f9";
		wait for Clk_period;
		Addr <=  "00000100110011";
		Trees_din <= x"0a03f104";
		wait for Clk_period;
		Addr <=  "00000100110100";
		Trees_din <= x"00a104f9";
		wait for Clk_period;
		Addr <=  "00000100110101";
		Trees_din <= x"ffca04f9";
		wait for Clk_period;
		Addr <=  "00000100110110";
		Trees_din <= x"061cb50c";
		wait for Clk_period;
		Addr <=  "00000100110111";
		Trees_din <= x"0515e908";
		wait for Clk_period;
		Addr <=  "00000100111000";
		Trees_din <= x"0113b304";
		wait for Clk_period;
		Addr <=  "00000100111001";
		Trees_din <= x"00b104f9";
		wait for Clk_period;
		Addr <=  "00000100111010";
		Trees_din <= x"007104f9";
		wait for Clk_period;
		Addr <=  "00000100111011";
		Trees_din <= x"fffc04f9";
		wait for Clk_period;
		Addr <=  "00000100111100";
		Trees_din <= x"ffa904f9";
		wait for Clk_period;
		Addr <=  "00000100111101";
		Trees_din <= x"ff7f04f9";
		wait for Clk_period;
		Addr <=  "00000100111110";
		Trees_din <= x"020b1e1c";
		wait for Clk_period;
		Addr <=  "00000100111111";
		Trees_din <= x"02030104";
		wait for Clk_period;
		Addr <=  "00000101000000";
		Trees_din <= x"ff64057d";
		wait for Clk_period;
		Addr <=  "00000101000001";
		Trees_din <= x"04007514";
		wait for Clk_period;
		Addr <=  "00000101000010";
		Trees_din <= x"05098d10";
		wait for Clk_period;
		Addr <=  "00000101000011";
		Trees_din <= x"000cbc08";
		wait for Clk_period;
		Addr <=  "00000101000100";
		Trees_din <= x"0a032304";
		wait for Clk_period;
		Addr <=  "00000101000101";
		Trees_din <= x"00ac057d";
		wait for Clk_period;
		Addr <=  "00000101000110";
		Trees_din <= x"ffb4057d";
		wait for Clk_period;
		Addr <=  "00000101000111";
		Trees_din <= x"11003904";
		wait for Clk_period;
		Addr <=  "00000101001000";
		Trees_din <= x"0045057d";
		wait for Clk_period;
		Addr <=  "00000101001001";
		Trees_din <= x"ff78057d";
		wait for Clk_period;
		Addr <=  "00000101001010";
		Trees_din <= x"ff75057d";
		wait for Clk_period;
		Addr <=  "00000101001011";
		Trees_din <= x"ff6c057d";
		wait for Clk_period;
		Addr <=  "00000101001100";
		Trees_din <= x"0113b318";
		wait for Clk_period;
		Addr <=  "00000101001101";
		Trees_din <= x"020f1914";
		wait for Clk_period;
		Addr <=  "00000101001110";
		Trees_din <= x"00f0ae08";
		wait for Clk_period;
		Addr <=  "00000101001111";
		Trees_din <= x"1100a704";
		wait for Clk_period;
		Addr <=  "00000101010000";
		Trees_din <= x"001e057d";
		wait for Clk_period;
		Addr <=  "00000101010001";
		Trees_din <= x"ff82057d";
		wait for Clk_period;
		Addr <=  "00000101010010";
		Trees_din <= x"06f98e04";
		wait for Clk_period;
		Addr <=  "00000101010011";
		Trees_din <= x"ff97057d";
		wait for Clk_period;
		Addr <=  "00000101010100";
		Trees_din <= x"0d03e704";
		wait for Clk_period;
		Addr <=  "00000101010101";
		Trees_din <= x"0094057d";
		wait for Clk_period;
		Addr <=  "00000101010110";
		Trees_din <= x"ffc7057d";
		wait for Clk_period;
		Addr <=  "00000101010111";
		Trees_din <= x"00a7057d";
		wait for Clk_period;
		Addr <=  "00000101011000";
		Trees_din <= x"021b0608";
		wait for Clk_period;
		Addr <=  "00000101011001";
		Trees_din <= x"02160e04";
		wait for Clk_period;
		Addr <=  "00000101011010";
		Trees_din <= x"ff6f057d";
		wait for Clk_period;
		Addr <=  "00000101011011";
		Trees_din <= x"fffd057d";
		wait for Clk_period;
		Addr <=  "00000101011100";
		Trees_din <= x"10fed404";
		wait for Clk_period;
		Addr <=  "00000101011101";
		Trees_din <= x"0017057d";
		wait for Clk_period;
		Addr <=  "00000101011110";
		Trees_din <= x"009f057d";
		wait for Clk_period;
		Addr <=  "00000101011111";
		Trees_din <= x"020b1e18";
		wait for Clk_period;
		Addr <=  "00000101100000";
		Trees_din <= x"02030104";
		wait for Clk_period;
		Addr <=  "00000101100001";
		Trees_din <= x"ff650601";
		wait for Clk_period;
		Addr <=  "00000101100010";
		Trees_din <= x"04009e10";
		wait for Clk_period;
		Addr <=  "00000101100011";
		Trees_din <= x"05098d0c";
		wait for Clk_period;
		Addr <=  "00000101100100";
		Trees_din <= x"000ec808";
		wait for Clk_period;
		Addr <=  "00000101100101";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00000101100110";
		Trees_din <= x"fff60601";
		wait for Clk_period;
		Addr <=  "00000101100111";
		Trees_din <= x"00b30601";
		wait for Clk_period;
		Addr <=  "00000101101000";
		Trees_din <= x"ff810601";
		wait for Clk_period;
		Addr <=  "00000101101001";
		Trees_din <= x"ff790601";
		wait for Clk_period;
		Addr <=  "00000101101010";
		Trees_din <= x"ff6c0601";
		wait for Clk_period;
		Addr <=  "00000101101011";
		Trees_din <= x"011fa028";
		wait for Clk_period;
		Addr <=  "00000101101100";
		Trees_din <= x"0210741c";
		wait for Clk_period;
		Addr <=  "00000101101101";
		Trees_din <= x"0402520c";
		wait for Clk_period;
		Addr <=  "00000101101110";
		Trees_din <= x"050ce108";
		wait for Clk_period;
		Addr <=  "00000101101111";
		Trees_din <= x"00f2af04";
		wait for Clk_period;
		Addr <=  "00000101110000";
		Trees_din <= x"00050601";
		wait for Clk_period;
		Addr <=  "00000101110001";
		Trees_din <= x"00970601";
		wait for Clk_period;
		Addr <=  "00000101110010";
		Trees_din <= x"ffa90601";
		wait for Clk_period;
		Addr <=  "00000101110011";
		Trees_din <= x"17004308";
		wait for Clk_period;
		Addr <=  "00000101110100";
		Trees_din <= x"04081e04";
		wait for Clk_period;
		Addr <=  "00000101110101";
		Trees_din <= x"00580601";
		wait for Clk_period;
		Addr <=  "00000101110110";
		Trees_din <= x"ff900601";
		wait for Clk_period;
		Addr <=  "00000101110111";
		Trees_din <= x"07005604";
		wait for Clk_period;
		Addr <=  "00000101111000";
		Trees_din <= x"fff70601";
		wait for Clk_period;
		Addr <=  "00000101111001";
		Trees_din <= x"ff5f0601";
		wait for Clk_period;
		Addr <=  "00000101111010";
		Trees_din <= x"0116f104";
		wait for Clk_period;
		Addr <=  "00000101111011";
		Trees_din <= x"00a30601";
		wait for Clk_period;
		Addr <=  "00000101111100";
		Trees_din <= x"13028804";
		wait for Clk_period;
		Addr <=  "00000101111101";
		Trees_din <= x"007d0601";
		wait for Clk_period;
		Addr <=  "00000101111110";
		Trees_din <= x"fffc0601";
		wait for Clk_period;
		Addr <=  "00000101111111";
		Trees_din <= x"ff8b0601";
		wait for Clk_period;
		Addr <=  "00000110000000";
		Trees_din <= x"020b1e28";
		wait for Clk_period;
		Addr <=  "00000110000001";
		Trees_din <= x"02030104";
		wait for Clk_period;
		Addr <=  "00000110000010";
		Trees_din <= x"ff6606b5";
		wait for Clk_period;
		Addr <=  "00000110000011";
		Trees_din <= x"04009e20";
		wait for Clk_period;
		Addr <=  "00000110000100";
		Trees_din <= x"07005810";
		wait for Clk_period;
		Addr <=  "00000110000101";
		Trees_din <= x"0c027f08";
		wait for Clk_period;
		Addr <=  "00000110000110";
		Trees_din <= x"06008804";
		wait for Clk_period;
		Addr <=  "00000110000111";
		Trees_din <= x"ff8306b5";
		wait for Clk_period;
		Addr <=  "00000110001000";
		Trees_din <= x"ffea06b5";
		wait for Clk_period;
		Addr <=  "00000110001001";
		Trees_din <= x"07005004";
		wait for Clk_period;
		Addr <=  "00000110001010";
		Trees_din <= x"005306b5";
		wait for Clk_period;
		Addr <=  "00000110001011";
		Trees_din <= x"ffad06b5";
		wait for Clk_period;
		Addr <=  "00000110001100";
		Trees_din <= x"1c003908";
		wait for Clk_period;
		Addr <=  "00000110001101";
		Trees_din <= x"05098d04";
		wait for Clk_period;
		Addr <=  "00000110001110";
		Trees_din <= x"00bd06b5";
		wait for Clk_period;
		Addr <=  "00000110001111";
		Trees_din <= x"ffb006b5";
		wait for Clk_period;
		Addr <=  "00000110010000";
		Trees_din <= x"02072404";
		wait for Clk_period;
		Addr <=  "00000110010001";
		Trees_din <= x"ff8c06b5";
		wait for Clk_period;
		Addr <=  "00000110010010";
		Trees_din <= x"002906b5";
		wait for Clk_period;
		Addr <=  "00000110010011";
		Trees_din <= x"ff6f06b5";
		wait for Clk_period;
		Addr <=  "00000110010100";
		Trees_din <= x"020f1920";
		wait for Clk_period;
		Addr <=  "00000110010101";
		Trees_din <= x"0402520c";
		wait for Clk_period;
		Addr <=  "00000110010110";
		Trees_din <= x"0506ce08";
		wait for Clk_period;
		Addr <=  "00000110010111";
		Trees_din <= x"07005b04";
		wait for Clk_period;
		Addr <=  "00000110011000";
		Trees_din <= x"009006b5";
		wait for Clk_period;
		Addr <=  "00000110011001";
		Trees_din <= x"fffe06b5";
		wait for Clk_period;
		Addr <=  "00000110011010";
		Trees_din <= x"fff806b5";
		wait for Clk_period;
		Addr <=  "00000110011011";
		Trees_din <= x"0700590c";
		wait for Clk_period;
		Addr <=  "00000110011100";
		Trees_din <= x"07005708";
		wait for Clk_period;
		Addr <=  "00000110011101";
		Trees_din <= x"00e76404";
		wait for Clk_period;
		Addr <=  "00000110011110";
		Trees_din <= x"ff9906b5";
		wait for Clk_period;
		Addr <=  "00000110011111";
		Trees_din <= x"006006b5";
		wait for Clk_period;
		Addr <=  "00000110100000";
		Trees_din <= x"ff4d06b5";
		wait for Clk_period;
		Addr <=  "00000110100001";
		Trees_din <= x"00eab204";
		wait for Clk_period;
		Addr <=  "00000110100010";
		Trees_din <= x"fff306b5";
		wait for Clk_period;
		Addr <=  "00000110100011";
		Trees_din <= x"005d06b5";
		wait for Clk_period;
		Addr <=  "00000110100100";
		Trees_din <= x"011fa010";
		wait for Clk_period;
		Addr <=  "00000110100101";
		Trees_din <= x"0515e90c";
		wait for Clk_period;
		Addr <=  "00000110100110";
		Trees_din <= x"0113b304";
		wait for Clk_period;
		Addr <=  "00000110100111";
		Trees_din <= x"00a006b5";
		wait for Clk_period;
		Addr <=  "00000110101000";
		Trees_din <= x"0213dd04";
		wait for Clk_period;
		Addr <=  "00000110101001";
		Trees_din <= x"ff9606b5";
		wait for Clk_period;
		Addr <=  "00000110101010";
		Trees_din <= x"008306b5";
		wait for Clk_period;
		Addr <=  "00000110101011";
		Trees_din <= x"fff806b5";
		wait for Clk_period;
		Addr <=  "00000110101100";
		Trees_din <= x"ffa006b5";
		wait for Clk_period;
		Addr <=  "00000110101101";
		Trees_din <= x"02083620";
		wait for Clk_period;
		Addr <=  "00000110101110";
		Trees_din <= x"02030104";
		wait for Clk_period;
		Addr <=  "00000110101111";
		Trees_din <= x"ff670759";
		wait for Clk_period;
		Addr <=  "00000110110000";
		Trees_din <= x"0a000f0c";
		wait for Clk_period;
		Addr <=  "00000110110001";
		Trees_din <= x"00067504";
		wait for Clk_period;
		Addr <=  "00000110110010";
		Trees_din <= x"ffac0759";
		wait for Clk_period;
		Addr <=  "00000110110011";
		Trees_din <= x"000cbc04";
		wait for Clk_period;
		Addr <=  "00000110110100";
		Trees_din <= x"00d40759";
		wait for Clk_period;
		Addr <=  "00000110110101";
		Trees_din <= x"ffae0759";
		wait for Clk_period;
		Addr <=  "00000110110110";
		Trees_din <= x"03fbf70c";
		wait for Clk_period;
		Addr <=  "00000110110111";
		Trees_din <= x"0c023808";
		wait for Clk_period;
		Addr <=  "00000110111000";
		Trees_din <= x"08005704";
		wait for Clk_period;
		Addr <=  "00000110111001";
		Trees_din <= x"ff930759";
		wait for Clk_period;
		Addr <=  "00000110111010";
		Trees_din <= x"fff30759";
		wait for Clk_period;
		Addr <=  "00000110111011";
		Trees_din <= x"00b00759";
		wait for Clk_period;
		Addr <=  "00000110111100";
		Trees_din <= x"ff6f0759";
		wait for Clk_period;
		Addr <=  "00000110111101";
		Trees_din <= x"020f1924";
		wait for Clk_period;
		Addr <=  "00000110111110";
		Trees_din <= x"00f1de08";
		wait for Clk_period;
		Addr <=  "00000110111111";
		Trees_din <= x"0ffe5204";
		wait for Clk_period;
		Addr <=  "00000111000000";
		Trees_din <= x"000b0759";
		wait for Clk_period;
		Addr <=  "00000111000001";
		Trees_din <= x"ff7b0759";
		wait for Clk_period;
		Addr <=  "00000111000010";
		Trees_din <= x"1700440c";
		wait for Clk_period;
		Addr <=  "00000111000011";
		Trees_din <= x"09055408";
		wait for Clk_period;
		Addr <=  "00000111000100";
		Trees_din <= x"0c002804";
		wait for Clk_period;
		Addr <=  "00000111000101";
		Trees_din <= x"00210759";
		wait for Clk_period;
		Addr <=  "00000111000110";
		Trees_din <= x"00870759";
		wait for Clk_period;
		Addr <=  "00000111000111";
		Trees_din <= x"ffee0759";
		wait for Clk_period;
		Addr <=  "00000111001000";
		Trees_din <= x"1401d808";
		wait for Clk_period;
		Addr <=  "00000111001001";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00000111001010";
		Trees_din <= x"ff670759";
		wait for Clk_period;
		Addr <=  "00000111001011";
		Trees_din <= x"00340759";
		wait for Clk_period;
		Addr <=  "00000111001100";
		Trees_din <= x"06fd9f04";
		wait for Clk_period;
		Addr <=  "00000111001101";
		Trees_din <= x"001c0759";
		wait for Clk_period;
		Addr <=  "00000111001110";
		Trees_din <= x"00660759";
		wait for Clk_period;
		Addr <=  "00000111001111";
		Trees_din <= x"011fa00c";
		wait for Clk_period;
		Addr <=  "00000111010000";
		Trees_din <= x"0113b304";
		wait for Clk_period;
		Addr <=  "00000111010001";
		Trees_din <= x"00990759";
		wait for Clk_period;
		Addr <=  "00000111010010";
		Trees_din <= x"0213dd04";
		wait for Clk_period;
		Addr <=  "00000111010011";
		Trees_din <= x"ff9f0759";
		wait for Clk_period;
		Addr <=  "00000111010100";
		Trees_din <= x"00800759";
		wait for Clk_period;
		Addr <=  "00000111010101";
		Trees_din <= x"ffa60759";
		wait for Clk_period;
		Addr <=  "00000111010110";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00000111010111";
		Trees_din <= x"02083624";
		wait for Clk_period;
		Addr <=  "00000111011000";
		Trees_din <= x"02030104";
		wait for Clk_period;
		Addr <=  "00000111011001";
		Trees_din <= x"ff6807f1";
		wait for Clk_period;
		Addr <=  "00000111011010";
		Trees_din <= x"0a000f10";
		wait for Clk_period;
		Addr <=  "00000111011011";
		Trees_din <= x"00067504";
		wait for Clk_period;
		Addr <=  "00000111011100";
		Trees_din <= x"ffb407f1";
		wait for Clk_period;
		Addr <=  "00000111011101";
		Trees_din <= x"1d00bd04";
		wait for Clk_period;
		Addr <=  "00000111011110";
		Trees_din <= x"fffd07f1";
		wait for Clk_period;
		Addr <=  "00000111011111";
		Trees_din <= x"1e006a04";
		wait for Clk_period;
		Addr <=  "00000111100000";
		Trees_din <= x"001f07f1";
		wait for Clk_period;
		Addr <=  "00000111100001";
		Trees_din <= x"00ba07f1";
		wait for Clk_period;
		Addr <=  "00000111100010";
		Trees_din <= x"03fbf70c";
		wait for Clk_period;
		Addr <=  "00000111100011";
		Trees_din <= x"06009f08";
		wait for Clk_period;
		Addr <=  "00000111100100";
		Trees_din <= x"08005804";
		wait for Clk_period;
		Addr <=  "00000111100101";
		Trees_din <= x"ff9b07f1";
		wait for Clk_period;
		Addr <=  "00000111100110";
		Trees_din <= x"ffee07f1";
		wait for Clk_period;
		Addr <=  "00000111100111";
		Trees_din <= x"00ab07f1";
		wait for Clk_period;
		Addr <=  "00000111101000";
		Trees_din <= x"ff7207f1";
		wait for Clk_period;
		Addr <=  "00000111101001";
		Trees_din <= x"020f1918";
		wait for Clk_period;
		Addr <=  "00000111101010";
		Trees_din <= x"00f1de08";
		wait for Clk_period;
		Addr <=  "00000111101011";
		Trees_din <= x"1f028804";
		wait for Clk_period;
		Addr <=  "00000111101100";
		Trees_din <= x"000507f1";
		wait for Clk_period;
		Addr <=  "00000111101101";
		Trees_din <= x"ff8107f1";
		wait for Clk_period;
		Addr <=  "00000111101110";
		Trees_din <= x"1402b50c";
		wait for Clk_period;
		Addr <=  "00000111101111";
		Trees_din <= x"04025208";
		wait for Clk_period;
		Addr <=  "00000111110000";
		Trees_din <= x"0c009604";
		wait for Clk_period;
		Addr <=  "00000111110001";
		Trees_din <= x"ffee07f1";
		wait for Clk_period;
		Addr <=  "00000111110010";
		Trees_din <= x"006807f1";
		wait for Clk_period;
		Addr <=  "00000111110011";
		Trees_din <= x"ff8a07f1";
		wait for Clk_period;
		Addr <=  "00000111110100";
		Trees_din <= x"007a07f1";
		wait for Clk_period;
		Addr <=  "00000111110101";
		Trees_din <= x"011fa00c";
		wait for Clk_period;
		Addr <=  "00000111110110";
		Trees_din <= x"0113b304";
		wait for Clk_period;
		Addr <=  "00000111110111";
		Trees_din <= x"009507f1";
		wait for Clk_period;
		Addr <=  "00000111111000";
		Trees_din <= x"0213dd04";
		wait for Clk_period;
		Addr <=  "00000111111001";
		Trees_din <= x"ffa607f1";
		wait for Clk_period;
		Addr <=  "00000111111010";
		Trees_din <= x"007707f1";
		wait for Clk_period;
		Addr <=  "00000111111011";
		Trees_din <= x"ffad07f1";
		wait for Clk_period;
		Addr <=  "00000111111100";
		Trees_din <= x"020b1e24";
		wait for Clk_period;
		Addr <=  "00000111111101";
		Trees_din <= x"02030104";
		wait for Clk_period;
		Addr <=  "00000111111110";
		Trees_din <= x"ff690895";
		wait for Clk_period;
		Addr <=  "00000111111111";
		Trees_din <= x"0400751c";
		wait for Clk_period;
		Addr <=  "00001000000000";
		Trees_din <= x"0700580c";
		wait for Clk_period;
		Addr <=  "00001000000001";
		Trees_din <= x"08004f08";
		wait for Clk_period;
		Addr <=  "00001000000010";
		Trees_din <= x"0c027704";
		wait for Clk_period;
		Addr <=  "00001000000011";
		Trees_din <= x"ffd40895";
		wait for Clk_period;
		Addr <=  "00001000000100";
		Trees_din <= x"00320895";
		wait for Clk_period;
		Addr <=  "00001000000101";
		Trees_din <= x"ff940895";
		wait for Clk_period;
		Addr <=  "00001000000110";
		Trees_din <= x"17004308";
		wait for Clk_period;
		Addr <=  "00001000000111";
		Trees_din <= x"17004204";
		wait for Clk_period;
		Addr <=  "00001000001000";
		Trees_din <= x"00210895";
		wait for Clk_period;
		Addr <=  "00001000001001";
		Trees_din <= x"00e40895";
		wait for Clk_period;
		Addr <=  "00001000001010";
		Trees_din <= x"02083604";
		wait for Clk_period;
		Addr <=  "00001000001011";
		Trees_din <= x"ffc20895";
		wait for Clk_period;
		Addr <=  "00001000001100";
		Trees_din <= x"002f0895";
		wait for Clk_period;
		Addr <=  "00001000001101";
		Trees_din <= x"ff7c0895";
		wait for Clk_period;
		Addr <=  "00001000001110";
		Trees_din <= x"0210741c";
		wait for Clk_period;
		Addr <=  "00001000001111";
		Trees_din <= x"00df9f04";
		wait for Clk_period;
		Addr <=  "00001000010000";
		Trees_din <= x"ff8d0895";
		wait for Clk_period;
		Addr <=  "00001000010001";
		Trees_din <= x"1a00490c";
		wait for Clk_period;
		Addr <=  "00001000010010";
		Trees_din <= x"00f95f08";
		wait for Clk_period;
		Addr <=  "00001000010011";
		Trees_din <= x"0efd3804";
		wait for Clk_period;
		Addr <=  "00001000010100";
		Trees_din <= x"004d0895";
		wait for Clk_period;
		Addr <=  "00001000010101";
		Trees_din <= x"ffd80895";
		wait for Clk_period;
		Addr <=  "00001000010110";
		Trees_din <= x"00810895";
		wait for Clk_period;
		Addr <=  "00001000010111";
		Trees_din <= x"0903c108";
		wait for Clk_period;
		Addr <=  "00001000011000";
		Trees_din <= x"0f013304";
		wait for Clk_period;
		Addr <=  "00001000011001";
		Trees_din <= x"ff780895";
		wait for Clk_period;
		Addr <=  "00001000011010";
		Trees_din <= x"00020895";
		wait for Clk_period;
		Addr <=  "00001000011011";
		Trees_din <= x"00480895";
		wait for Clk_period;
		Addr <=  "00001000011100";
		Trees_din <= x"0412100c";
		wait for Clk_period;
		Addr <=  "00001000011101";
		Trees_din <= x"02128c08";
		wait for Clk_period;
		Addr <=  "00001000011110";
		Trees_din <= x"00e88e04";
		wait for Clk_period;
		Addr <=  "00001000011111";
		Trees_din <= x"ffda0895";
		wait for Clk_period;
		Addr <=  "00001000100000";
		Trees_din <= x"00820895";
		wait for Clk_period;
		Addr <=  "00001000100001";
		Trees_din <= x"00960895";
		wait for Clk_period;
		Addr <=  "00001000100010";
		Trees_din <= x"021ddb04";
		wait for Clk_period;
		Addr <=  "00001000100011";
		Trees_din <= x"ffad0895";
		wait for Clk_period;
		Addr <=  "00001000100100";
		Trees_din <= x"00620895";
		wait for Clk_period;
		Addr <=  "00001000100101";
		Trees_din <= x"02083620";
		wait for Clk_period;
		Addr <=  "00001000100110";
		Trees_din <= x"02030104";
		wait for Clk_period;
		Addr <=  "00001000100111";
		Trees_din <= x"ff6a0931";
		wait for Clk_period;
		Addr <=  "00001000101000";
		Trees_din <= x"13028710";
		wait for Clk_period;
		Addr <=  "00001000101001";
		Trees_din <= x"03fbeb0c";
		wait for Clk_period;
		Addr <=  "00001000101010";
		Trees_din <= x"06feb104";
		wait for Clk_period;
		Addr <=  "00001000101011";
		Trees_din <= x"ffa90931";
		wait for Clk_period;
		Addr <=  "00001000101100";
		Trees_din <= x"09043804";
		wait for Clk_period;
		Addr <=  "00001000101101";
		Trees_din <= x"ffff0931";
		wait for Clk_period;
		Addr <=  "00001000101110";
		Trees_din <= x"00590931";
		wait for Clk_period;
		Addr <=  "00001000101111";
		Trees_din <= x"ff7a0931";
		wait for Clk_period;
		Addr <=  "00001000110000";
		Trees_din <= x"01fcd508";
		wait for Clk_period;
		Addr <=  "00001000110001";
		Trees_din <= x"10012e04";
		wait for Clk_period;
		Addr <=  "00001000110010";
		Trees_din <= x"fff60931";
		wait for Clk_period;
		Addr <=  "00001000110011";
		Trees_din <= x"00d80931";
		wait for Clk_period;
		Addr <=  "00001000110100";
		Trees_din <= x"ffa30931";
		wait for Clk_period;
		Addr <=  "00001000110101";
		Trees_din <= x"02107420";
		wait for Clk_period;
		Addr <=  "00001000110110";
		Trees_din <= x"00f2af08";
		wait for Clk_period;
		Addr <=  "00001000110111";
		Trees_din <= x"10fe2904";
		wait for Clk_period;
		Addr <=  "00001000111000";
		Trees_din <= x"00170931";
		wait for Clk_period;
		Addr <=  "00001000111001";
		Trees_din <= x"ff8d0931";
		wait for Clk_period;
		Addr <=  "00001000111010";
		Trees_din <= x"1700440c";
		wait for Clk_period;
		Addr <=  "00001000111011";
		Trees_din <= x"09055408";
		wait for Clk_period;
		Addr <=  "00001000111100";
		Trees_din <= x"0c005104";
		wait for Clk_period;
		Addr <=  "00001000111101";
		Trees_din <= x"001b0931";
		wait for Clk_period;
		Addr <=  "00001000111110";
		Trees_din <= x"00790931";
		wait for Clk_period;
		Addr <=  "00001000111111";
		Trees_din <= x"fffd0931";
		wait for Clk_period;
		Addr <=  "00001001000000";
		Trees_din <= x"0fff2e04";
		wait for Clk_period;
		Addr <=  "00001001000001";
		Trees_din <= x"ff9e0931";
		wait for Clk_period;
		Addr <=  "00001001000010";
		Trees_din <= x"04007504";
		wait for Clk_period;
		Addr <=  "00001001000011";
		Trees_din <= x"005d0931";
		wait for Clk_period;
		Addr <=  "00001001000100";
		Trees_din <= x"ffe30931";
		wait for Clk_period;
		Addr <=  "00001001000101";
		Trees_din <= x"0412100c";
		wait for Clk_period;
		Addr <=  "00001001000110";
		Trees_din <= x"02117808";
		wait for Clk_period;
		Addr <=  "00001001000111";
		Trees_din <= x"03fe0b04";
		wait for Clk_period;
		Addr <=  "00001001001000";
		Trees_din <= x"005d0931";
		wait for Clk_period;
		Addr <=  "00001001001001";
		Trees_din <= x"ffff0931";
		wait for Clk_period;
		Addr <=  "00001001001010";
		Trees_din <= x"00900931";
		wait for Clk_period;
		Addr <=  "00001001001011";
		Trees_din <= x"00110931";
		wait for Clk_period;
		Addr <=  "00001001001100";
		Trees_din <= x"020b1e24";
		wait for Clk_period;
		Addr <=  "00001001001101";
		Trees_din <= x"02030104";
		wait for Clk_period;
		Addr <=  "00001001001110";
		Trees_din <= x"ff6b09c5";
		wait for Clk_period;
		Addr <=  "00001001001111";
		Trees_din <= x"07005808";
		wait for Clk_period;
		Addr <=  "00001001010000";
		Trees_din <= x"04fd2604";
		wait for Clk_period;
		Addr <=  "00001001010001";
		Trees_din <= x"000609c5";
		wait for Clk_period;
		Addr <=  "00001001010010";
		Trees_din <= x"ff9109c5";
		wait for Clk_period;
		Addr <=  "00001001010011";
		Trees_din <= x"03fbf70c";
		wait for Clk_period;
		Addr <=  "00001001010100";
		Trees_din <= x"03fbd808";
		wait for Clk_period;
		Addr <=  "00001001010101";
		Trees_din <= x"14028e04";
		wait for Clk_period;
		Addr <=  "00001001010110";
		Trees_din <= x"ffd809c5";
		wait for Clk_period;
		Addr <=  "00001001010111";
		Trees_din <= x"004309c5";
		wait for Clk_period;
		Addr <=  "00001001011000";
		Trees_din <= x"00e109c5";
		wait for Clk_period;
		Addr <=  "00001001011001";
		Trees_din <= x"0a000104";
		wait for Clk_period;
		Addr <=  "00001001011010";
		Trees_din <= x"004809c5";
		wait for Clk_period;
		Addr <=  "00001001011011";
		Trees_din <= x"02088f04";
		wait for Clk_period;
		Addr <=  "00001001011100";
		Trees_din <= x"ff9009c5";
		wait for Clk_period;
		Addr <=  "00001001011101";
		Trees_din <= x"000a09c5";
		wait for Clk_period;
		Addr <=  "00001001011110";
		Trees_din <= x"02107418";
		wait for Clk_period;
		Addr <=  "00001001011111";
		Trees_din <= x"0402520c";
		wait for Clk_period;
		Addr <=  "00001001100000";
		Trees_din <= x"0c007308";
		wait for Clk_period;
		Addr <=  "00001001100001";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00001001100010";
		Trees_din <= x"003e09c5";
		wait for Clk_period;
		Addr <=  "00001001100011";
		Trees_din <= x"ffee09c5";
		wait for Clk_period;
		Addr <=  "00001001100100";
		Trees_din <= x"007009c5";
		wait for Clk_period;
		Addr <=  "00001001100101";
		Trees_din <= x"07005908";
		wait for Clk_period;
		Addr <=  "00001001100110";
		Trees_din <= x"07005504";
		wait for Clk_period;
		Addr <=  "00001001100111";
		Trees_din <= x"000a09c5";
		wait for Clk_period;
		Addr <=  "00001001101000";
		Trees_din <= x"ff7c09c5";
		wait for Clk_period;
		Addr <=  "00001001101001";
		Trees_din <= x"003009c5";
		wait for Clk_period;
		Addr <=  "00001001101010";
		Trees_din <= x"0412100c";
		wait for Clk_period;
		Addr <=  "00001001101011";
		Trees_din <= x"02128c08";
		wait for Clk_period;
		Addr <=  "00001001101100";
		Trees_din <= x"00e88e04";
		wait for Clk_period;
		Addr <=  "00001001101101";
		Trees_din <= x"ffdc09c5";
		wait for Clk_period;
		Addr <=  "00001001101110";
		Trees_din <= x"007609c5";
		wait for Clk_period;
		Addr <=  "00001001101111";
		Trees_din <= x"008f09c5";
		wait for Clk_period;
		Addr <=  "00001001110000";
		Trees_din <= x"000d09c5";
		wait for Clk_period;
		Addr <=  "00001001110001";
		Trees_din <= x"02030104";
		wait for Clk_period;
		Addr <=  "00001001110010";
		Trees_din <= x"ff6d0a39";
		wait for Clk_period;
		Addr <=  "00001001110011";
		Trees_din <= x"020f1924";
		wait for Clk_period;
		Addr <=  "00001001110100";
		Trees_din <= x"00f95f08";
		wait for Clk_period;
		Addr <=  "00001001110101";
		Trees_din <= x"0ef8cc04";
		wait for Clk_period;
		Addr <=  "00001001110110";
		Trees_din <= x"00100a39";
		wait for Clk_period;
		Addr <=  "00001001110111";
		Trees_din <= x"ff8a0a39";
		wait for Clk_period;
		Addr <=  "00001001111000";
		Trees_din <= x"03fbf710";
		wait for Clk_period;
		Addr <=  "00001001111001";
		Trees_din <= x"1401a608";
		wait for Clk_period;
		Addr <=  "00001001111010";
		Trees_din <= x"03fac204";
		wait for Clk_period;
		Addr <=  "00001001111011";
		Trees_din <= x"00380a39";
		wait for Clk_period;
		Addr <=  "00001001111100";
		Trees_din <= x"ffb70a39";
		wait for Clk_period;
		Addr <=  "00001001111101";
		Trees_din <= x"06fe2704";
		wait for Clk_period;
		Addr <=  "00001001111110";
		Trees_din <= x"00230a39";
		wait for Clk_period;
		Addr <=  "00001001111111";
		Trees_din <= x"00b30a39";
		wait for Clk_period;
		Addr <=  "00001010000000";
		Trees_din <= x"0a000104";
		wait for Clk_period;
		Addr <=  "00001010000001";
		Trees_din <= x"00440a39";
		wait for Clk_period;
		Addr <=  "00001010000010";
		Trees_din <= x"02088f04";
		wait for Clk_period;
		Addr <=  "00001010000011";
		Trees_din <= x"ff890a39";
		wait for Clk_period;
		Addr <=  "00001010000100";
		Trees_din <= x"000b0a39";
		wait for Clk_period;
		Addr <=  "00001010000101";
		Trees_din <= x"00c0270c";
		wait for Clk_period;
		Addr <=  "00001010000110";
		Trees_din <= x"021b0604";
		wait for Clk_period;
		Addr <=  "00001010000111";
		Trees_din <= x"ffb20a39";
		wait for Clk_period;
		Addr <=  "00001010001000";
		Trees_din <= x"0f007904";
		wait for Clk_period;
		Addr <=  "00001010001001";
		Trees_din <= x"00130a39";
		wait for Clk_period;
		Addr <=  "00001010001010";
		Trees_din <= x"007c0a39";
		wait for Clk_period;
		Addr <=  "00001010001011";
		Trees_din <= x"18004e04";
		wait for Clk_period;
		Addr <=  "00001010001100";
		Trees_din <= x"008c0a39";
		wait for Clk_period;
		Addr <=  "00001010001101";
		Trees_din <= x"00280a39";
		wait for Clk_period;
		Addr <=  "00001010001110";
		Trees_din <= x"02030104";
		wait for Clk_period;
		Addr <=  "00001010001111";
		Trees_din <= x"ff6f0aad";
		wait for Clk_period;
		Addr <=  "00001010010000";
		Trees_din <= x"020f1928";
		wait for Clk_period;
		Addr <=  "00001010010001";
		Trees_din <= x"04007518";
		wait for Clk_period;
		Addr <=  "00001010010010";
		Trees_din <= x"0506ce10";
		wait for Clk_period;
		Addr <=  "00001010010011";
		Trees_din <= x"03fbf708";
		wait for Clk_period;
		Addr <=  "00001010010100";
		Trees_din <= x"17003f04";
		wait for Clk_period;
		Addr <=  "00001010010101";
		Trees_din <= x"00070aad";
		wait for Clk_period;
		Addr <=  "00001010010110";
		Trees_din <= x"00990aad";
		wait for Clk_period;
		Addr <=  "00001010010111";
		Trees_din <= x"000cbc04";
		wait for Clk_period;
		Addr <=  "00001010011000";
		Trees_din <= x"00320aad";
		wait for Clk_period;
		Addr <=  "00001010011001";
		Trees_din <= x"ffb10aad";
		wait for Clk_period;
		Addr <=  "00001010011010";
		Trees_din <= x"02088f04";
		wait for Clk_period;
		Addr <=  "00001010011011";
		Trees_din <= x"ffa20aad";
		wait for Clk_period;
		Addr <=  "00001010011100";
		Trees_din <= x"00010aad";
		wait for Clk_period;
		Addr <=  "00001010011101";
		Trees_din <= x"08005a0c";
		wait for Clk_period;
		Addr <=  "00001010011110";
		Trees_din <= x"06fdd508";
		wait for Clk_period;
		Addr <=  "00001010011111";
		Trees_din <= x"1402bc04";
		wait for Clk_period;
		Addr <=  "00001010100000";
		Trees_din <= x"ffc30aad";
		wait for Clk_period;
		Addr <=  "00001010100001";
		Trees_din <= x"00240aad";
		wait for Clk_period;
		Addr <=  "00001010100010";
		Trees_din <= x"ff8f0aad";
		wait for Clk_period;
		Addr <=  "00001010100011";
		Trees_din <= x"001d0aad";
		wait for Clk_period;
		Addr <=  "00001010100100";
		Trees_din <= x"011a8c0c";
		wait for Clk_period;
		Addr <=  "00001010100101";
		Trees_din <= x"02117808";
		wait for Clk_period;
		Addr <=  "00001010100110";
		Trees_din <= x"06030404";
		wait for Clk_period;
		Addr <=  "00001010100111";
		Trees_din <= x"005f0aad";
		wait for Clk_period;
		Addr <=  "00001010101000";
		Trees_din <= x"ffec0aad";
		wait for Clk_period;
		Addr <=  "00001010101001";
		Trees_din <= x"00880aad";
		wait for Clk_period;
		Addr <=  "00001010101010";
		Trees_din <= x"ffec0aad";
		wait for Clk_period;
		Addr <=  "00001010101011";
		Trees_din <= x"02030104";
		wait for Clk_period;
		Addr <=  "00001010101100";
		Trees_din <= x"ff710b21";
		wait for Clk_period;
		Addr <=  "00001010101101";
		Trees_din <= x"020f1928";
		wait for Clk_period;
		Addr <=  "00001010101110";
		Trees_din <= x"04007518";
		wait for Clk_period;
		Addr <=  "00001010101111";
		Trees_din <= x"05058710";
		wait for Clk_period;
		Addr <=  "00001010110000";
		Trees_din <= x"07005808";
		wait for Clk_period;
		Addr <=  "00001010110001";
		Trees_din <= x"02072404";
		wait for Clk_period;
		Addr <=  "00001010110010";
		Trees_din <= x"ffc50b21";
		wait for Clk_period;
		Addr <=  "00001010110011";
		Trees_din <= x"003e0b21";
		wait for Clk_period;
		Addr <=  "00001010110100";
		Trees_din <= x"1d00ba04";
		wait for Clk_period;
		Addr <=  "00001010110101";
		Trees_din <= x"00050b21";
		wait for Clk_period;
		Addr <=  "00001010110110";
		Trees_din <= x"008f0b21";
		wait for Clk_period;
		Addr <=  "00001010110111";
		Trees_din <= x"07005a04";
		wait for Clk_period;
		Addr <=  "00001010111000";
		Trees_din <= x"ffb20b21";
		wait for Clk_period;
		Addr <=  "00001010111001";
		Trees_din <= x"001a0b21";
		wait for Clk_period;
		Addr <=  "00001010111010";
		Trees_din <= x"08005a0c";
		wait for Clk_period;
		Addr <=  "00001010111011";
		Trees_din <= x"06fdd508";
		wait for Clk_period;
		Addr <=  "00001010111100";
		Trees_din <= x"10011f04";
		wait for Clk_period;
		Addr <=  "00001010111101";
		Trees_din <= x"ffd30b21";
		wait for Clk_period;
		Addr <=  "00001010111110";
		Trees_din <= x"00130b21";
		wait for Clk_period;
		Addr <=  "00001010111111";
		Trees_din <= x"ff960b21";
		wait for Clk_period;
		Addr <=  "00001011000000";
		Trees_din <= x"00190b21";
		wait for Clk_period;
		Addr <=  "00001011000001";
		Trees_din <= x"00c0270c";
		wait for Clk_period;
		Addr <=  "00001011000010";
		Trees_din <= x"021ddb08";
		wait for Clk_period;
		Addr <=  "00001011000011";
		Trees_din <= x"0217b304";
		wait for Clk_period;
		Addr <=  "00001011000100";
		Trees_din <= x"ffad0b21";
		wait for Clk_period;
		Addr <=  "00001011000101";
		Trees_din <= x"fffe0b21";
		wait for Clk_period;
		Addr <=  "00001011000110";
		Trees_din <= x"00720b21";
		wait for Clk_period;
		Addr <=  "00001011000111";
		Trees_din <= x"00800b21";
		wait for Clk_period;
		Addr <=  "00001011001000";
		Trees_din <= x"02030104";
		wait for Clk_period;
		Addr <=  "00001011001001";
		Trees_din <= x"ff740b7d";
		wait for Clk_period;
		Addr <=  "00001011001010";
		Trees_din <= x"02107420";
		wait for Clk_period;
		Addr <=  "00001011001011";
		Trees_din <= x"00f95f08";
		wait for Clk_period;
		Addr <=  "00001011001100";
		Trees_din <= x"0fff3804";
		wait for Clk_period;
		Addr <=  "00001011001101";
		Trees_din <= x"fffb0b7d";
		wait for Clk_period;
		Addr <=  "00001011001110";
		Trees_din <= x"ffa10b7d";
		wait for Clk_period;
		Addr <=  "00001011001111";
		Trees_din <= x"1700440c";
		wait for Clk_period;
		Addr <=  "00001011010000";
		Trees_din <= x"17004208";
		wait for Clk_period;
		Addr <=  "00001011010001";
		Trees_din <= x"02088f04";
		wait for Clk_period;
		Addr <=  "00001011010010";
		Trees_din <= x"ffc70b7d";
		wait for Clk_period;
		Addr <=  "00001011010011";
		Trees_din <= x"00480b7d";
		wait for Clk_period;
		Addr <=  "00001011010100";
		Trees_din <= x"008b0b7d";
		wait for Clk_period;
		Addr <=  "00001011010101";
		Trees_din <= x"07005a08";
		wait for Clk_period;
		Addr <=  "00001011010110";
		Trees_din <= x"14016204";
		wait for Clk_period;
		Addr <=  "00001011010111";
		Trees_din <= x"ff9f0b7d";
		wait for Clk_period;
		Addr <=  "00001011011000";
		Trees_din <= x"ffee0b7d";
		wait for Clk_period;
		Addr <=  "00001011011001";
		Trees_din <= x"00170b7d";
		wait for Clk_period;
		Addr <=  "00001011011010";
		Trees_din <= x"04121008";
		wait for Clk_period;
		Addr <=  "00001011011011";
		Trees_din <= x"02128c04";
		wait for Clk_period;
		Addr <=  "00001011011100";
		Trees_din <= x"002e0b7d";
		wait for Clk_period;
		Addr <=  "00001011011101";
		Trees_din <= x"00810b7d";
		wait for Clk_period;
		Addr <=  "00001011011110";
		Trees_din <= x"00020b7d";
		wait for Clk_period;
		Addr <=  "00001011011111";
		Trees_din <= x"02030104";
		wait for Clk_period;
		Addr <=  "00001011100000";
		Trees_din <= x"ff780be1";
		wait for Clk_period;
		Addr <=  "00001011100001";
		Trees_din <= x"020f1920";
		wait for Clk_period;
		Addr <=  "00001011100010";
		Trees_din <= x"1200940c";
		wait for Clk_period;
		Addr <=  "00001011100011";
		Trees_din <= x"03fb8804";
		wait for Clk_period;
		Addr <=  "00001011100100";
		Trees_din <= x"000f0be1";
		wait for Clk_period;
		Addr <=  "00001011100101";
		Trees_din <= x"01fdf904";
		wait for Clk_period;
		Addr <=  "00001011100110";
		Trees_din <= x"ffdd0be1";
		wait for Clk_period;
		Addr <=  "00001011100111";
		Trees_din <= x"ff980be1";
		wait for Clk_period;
		Addr <=  "00001011101000";
		Trees_din <= x"13027f0c";
		wait for Clk_period;
		Addr <=  "00001011101001";
		Trees_din <= x"020bd208";
		wait for Clk_period;
		Addr <=  "00001011101010";
		Trees_din <= x"13fae004";
		wait for Clk_period;
		Addr <=  "00001011101011";
		Trees_din <= x"00070be1";
		wait for Clk_period;
		Addr <=  "00001011101100";
		Trees_din <= x"ffa80be1";
		wait for Clk_period;
		Addr <=  "00001011101101";
		Trees_din <= x"002f0be1";
		wait for Clk_period;
		Addr <=  "00001011101110";
		Trees_din <= x"17003e04";
		wait for Clk_period;
		Addr <=  "00001011101111";
		Trees_din <= x"00030be1";
		wait for Clk_period;
		Addr <=  "00001011110000";
		Trees_din <= x"00830be1";
		wait for Clk_period;
		Addr <=  "00001011110001";
		Trees_din <= x"0113b308";
		wait for Clk_period;
		Addr <=  "00001011110010";
		Trees_din <= x"05098d04";
		wait for Clk_period;
		Addr <=  "00001011110011";
		Trees_din <= x"00800be1";
		wait for Clk_period;
		Addr <=  "00001011110100";
		Trees_din <= x"001e0be1";
		wait for Clk_period;
		Addr <=  "00001011110101";
		Trees_din <= x"021ddb04";
		wait for Clk_period;
		Addr <=  "00001011110110";
		Trees_din <= x"ffbe0be1";
		wait for Clk_period;
		Addr <=  "00001011110111";
		Trees_din <= x"00510be1";
		wait for Clk_period;
		Addr <=  "00001011111000";
		Trees_din <= x"02030104";
		wait for Clk_period;
		Addr <=  "00001011111001";
		Trees_din <= x"ff7c0c3d";
		wait for Clk_period;
		Addr <=  "00001011111010";
		Trees_din <= x"02117824";
		wait for Clk_period;
		Addr <=  "00001011111011";
		Trees_din <= x"04025218";
		wait for Clk_period;
		Addr <=  "00001011111100";
		Trees_din <= x"0506f710";
		wait for Clk_period;
		Addr <=  "00001011111101";
		Trees_din <= x"03fbf708";
		wait for Clk_period;
		Addr <=  "00001011111110";
		Trees_din <= x"12009a04";
		wait for Clk_period;
		Addr <=  "00001011111111";
		Trees_din <= x"007b0c3d";
		wait for Clk_period;
		Addr <=  "00001100000000";
		Trees_din <= x"00110c3d";
		wait for Clk_period;
		Addr <=  "00001100000001";
		Trees_din <= x"13011b04";
		wait for Clk_period;
		Addr <=  "00001100000010";
		Trees_din <= x"ffdf0c3d";
		wait for Clk_period;
		Addr <=  "00001100000011";
		Trees_din <= x"00280c3d";
		wait for Clk_period;
		Addr <=  "00001100000100";
		Trees_din <= x"0c016d04";
		wait for Clk_period;
		Addr <=  "00001100000101";
		Trees_din <= x"ffb40c3d";
		wait for Clk_period;
		Addr <=  "00001100000110";
		Trees_din <= x"00040c3d";
		wait for Clk_period;
		Addr <=  "00001100000111";
		Trees_din <= x"07005908";
		wait for Clk_period;
		Addr <=  "00001100001000";
		Trees_din <= x"07005504";
		wait for Clk_period;
		Addr <=  "00001100001001";
		Trees_din <= x"fff40c3d";
		wait for Clk_period;
		Addr <=  "00001100001010";
		Trees_din <= x"ff980c3d";
		wait for Clk_period;
		Addr <=  "00001100001011";
		Trees_din <= x"000a0c3d";
		wait for Clk_period;
		Addr <=  "00001100001100";
		Trees_din <= x"0410ae04";
		wait for Clk_period;
		Addr <=  "00001100001101";
		Trees_din <= x"00740c3d";
		wait for Clk_period;
		Addr <=  "00001100001110";
		Trees_din <= x"000c0c3d";
		wait for Clk_period;
		Addr <=  "00001100001111";
		Trees_din <= x"020b1e18";
		wait for Clk_period;
		Addr <=  "00001100010000";
		Trees_din <= x"02030104";
		wait for Clk_period;
		Addr <=  "00001100010001";
		Trees_din <= x"ff810ca1";
		wait for Clk_period;
		Addr <=  "00001100010010";
		Trees_din <= x"07005908";
		wait for Clk_period;
		Addr <=  "00001100010011";
		Trees_din <= x"0a000f04";
		wait for Clk_period;
		Addr <=  "00001100010100";
		Trees_din <= x"000a0ca1";
		wait for Clk_period;
		Addr <=  "00001100010101";
		Trees_din <= x"ff9f0ca1";
		wait for Clk_period;
		Addr <=  "00001100010110";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00001100010111";
		Trees_din <= x"00650ca1";
		wait for Clk_period;
		Addr <=  "00001100011000";
		Trees_din <= x"14031104";
		wait for Clk_period;
		Addr <=  "00001100011001";
		Trees_din <= x"ffcd0ca1";
		wait for Clk_period;
		Addr <=  "00001100011010";
		Trees_din <= x"00110ca1";
		wait for Clk_period;
		Addr <=  "00001100011011";
		Trees_din <= x"0113b314";
		wait for Clk_period;
		Addr <=  "00001100011100";
		Trees_din <= x"020fd90c";
		wait for Clk_period;
		Addr <=  "00001100011101";
		Trees_din <= x"1a004908";
		wait for Clk_period;
		Addr <=  "00001100011110";
		Trees_din <= x"00f95f04";
		wait for Clk_period;
		Addr <=  "00001100011111";
		Trees_din <= x"fffb0ca1";
		wait for Clk_period;
		Addr <=  "00001100100000";
		Trees_din <= x"00560ca1";
		wait for Clk_period;
		Addr <=  "00001100100001";
		Trees_din <= x"ffda0ca1";
		wait for Clk_period;
		Addr <=  "00001100100010";
		Trees_din <= x"05098d04";
		wait for Clk_period;
		Addr <=  "00001100100011";
		Trees_din <= x"007a0ca1";
		wait for Clk_period;
		Addr <=  "00001100100100";
		Trees_din <= x"001d0ca1";
		wait for Clk_period;
		Addr <=  "00001100100101";
		Trees_din <= x"13fce404";
		wait for Clk_period;
		Addr <=  "00001100100110";
		Trees_din <= x"001c0ca1";
		wait for Clk_period;
		Addr <=  "00001100100111";
		Trees_din <= x"ffda0ca1";
		wait for Clk_period;
		Addr <=  "00001100101000";
		Trees_din <= x"020b1e18";
		wait for Clk_period;
		Addr <=  "00001100101001";
		Trees_din <= x"02030104";
		wait for Clk_period;
		Addr <=  "00001100101010";
		Trees_din <= x"ff860cfd";
		wait for Clk_period;
		Addr <=  "00001100101011";
		Trees_din <= x"1302870c";
		wait for Clk_period;
		Addr <=  "00001100101100";
		Trees_din <= x"02072404";
		wait for Clk_period;
		Addr <=  "00001100101101";
		Trees_din <= x"ffad0cfd";
		wait for Clk_period;
		Addr <=  "00001100101110";
		Trees_din <= x"07005704";
		wait for Clk_period;
		Addr <=  "00001100101111";
		Trees_din <= x"ffdf0cfd";
		wait for Clk_period;
		Addr <=  "00001100110000";
		Trees_din <= x"000d0cfd";
		wait for Clk_period;
		Addr <=  "00001100110001";
		Trees_din <= x"1b00f604";
		wait for Clk_period;
		Addr <=  "00001100110010";
		Trees_din <= x"00570cfd";
		wait for Clk_period;
		Addr <=  "00001100110011";
		Trees_din <= x"ffe20cfd";
		wait for Clk_period;
		Addr <=  "00001100110100";
		Trees_din <= x"02128c10";
		wait for Clk_period;
		Addr <=  "00001100110101";
		Trees_din <= x"00df9f04";
		wait for Clk_period;
		Addr <=  "00001100110110";
		Trees_din <= x"ffb10cfd";
		wait for Clk_period;
		Addr <=  "00001100110111";
		Trees_din <= x"08005604";
		wait for Clk_period;
		Addr <=  "00001100111000";
		Trees_din <= x"00550cfd";
		wait for Clk_period;
		Addr <=  "00001100111001";
		Trees_din <= x"09fcb804";
		wait for Clk_period;
		Addr <=  "00001100111010";
		Trees_din <= x"ffce0cfd";
		wait for Clk_period;
		Addr <=  "00001100111011";
		Trees_din <= x"003a0cfd";
		wait for Clk_period;
		Addr <=  "00001100111100";
		Trees_din <= x"04121004";
		wait for Clk_period;
		Addr <=  "00001100111101";
		Trees_din <= x"00700cfd";
		wait for Clk_period;
		Addr <=  "00001100111110";
		Trees_din <= x"000a0cfd";
		wait for Clk_period;
		Addr <=  "00001100111111";
		Trees_din <= x"020b1e14";
		wait for Clk_period;
		Addr <=  "00001101000000";
		Trees_din <= x"03fbf708";
		wait for Clk_period;
		Addr <=  "00001101000001";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00001101000010";
		Trees_din <= x"ffcd0d49";
		wait for Clk_period;
		Addr <=  "00001101000011";
		Trees_din <= x"00380d49";
		wait for Clk_period;
		Addr <=  "00001101000100";
		Trees_din <= x"0a000104";
		wait for Clk_period;
		Addr <=  "00001101000101";
		Trees_din <= x"000f0d49";
		wait for Clk_period;
		Addr <=  "00001101000110";
		Trees_din <= x"02088f04";
		wait for Clk_period;
		Addr <=  "00001101000111";
		Trees_din <= x"ff820d49";
		wait for Clk_period;
		Addr <=  "00001101001000";
		Trees_din <= x"fff20d49";
		wait for Clk_period;
		Addr <=  "00001101001001";
		Trees_din <= x"02128c0c";
		wait for Clk_period;
		Addr <=  "00001101001010";
		Trees_din <= x"00df9f04";
		wait for Clk_period;
		Addr <=  "00001101001011";
		Trees_din <= x"ffb70d49";
		wait for Clk_period;
		Addr <=  "00001101001100";
		Trees_din <= x"1a004904";
		wait for Clk_period;
		Addr <=  "00001101001101";
		Trees_din <= x"00490d49";
		wait for Clk_period;
		Addr <=  "00001101001110";
		Trees_din <= x"fff90d49";
		wait for Clk_period;
		Addr <=  "00001101001111";
		Trees_din <= x"0fff0604";
		wait for Clk_period;
		Addr <=  "00001101010000";
		Trees_din <= x"00170d49";
		wait for Clk_period;
		Addr <=  "00001101010001";
		Trees_din <= x"00670d49";
		wait for Clk_period;
		Addr <=  "00001101010010";
		Trees_din <= x"020b1e14";
		wait for Clk_period;
		Addr <=  "00001101010011";
		Trees_din <= x"02030104";
		wait for Clk_period;
		Addr <=  "00001101010100";
		Trees_din <= x"ff900d95";
		wait for Clk_period;
		Addr <=  "00001101010101";
		Trees_din <= x"00071308";
		wait for Clk_period;
		Addr <=  "00001101010110";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00001101010111";
		Trees_din <= x"ffae0d95";
		wait for Clk_period;
		Addr <=  "00001101011000";
		Trees_din <= x"fff70d95";
		wait for Clk_period;
		Addr <=  "00001101011001";
		Trees_din <= x"13028704";
		wait for Clk_period;
		Addr <=  "00001101011010";
		Trees_din <= x"ffe70d95";
		wait for Clk_period;
		Addr <=  "00001101011011";
		Trees_din <= x"004c0d95";
		wait for Clk_period;
		Addr <=  "00001101011100";
		Trees_din <= x"02159b10";
		wait for Clk_period;
		Addr <=  "00001101011101";
		Trees_din <= x"00df9f04";
		wait for Clk_period;
		Addr <=  "00001101011110";
		Trees_din <= x"ffb50d95";
		wait for Clk_period;
		Addr <=  "00001101011111";
		Trees_din <= x"08005604";
		wait for Clk_period;
		Addr <=  "00001101100000";
		Trees_din <= x"00520d95";
		wait for Clk_period;
		Addr <=  "00001101100001";
		Trees_din <= x"09fcb804";
		wait for Clk_period;
		Addr <=  "00001101100010";
		Trees_din <= x"ffd80d95";
		wait for Clk_period;
		Addr <=  "00001101100011";
		Trees_din <= x"00380d95";
		wait for Clk_period;
		Addr <=  "00001101100100";
		Trees_din <= x"005e0d95";
		wait for Clk_period;
		Addr <=  "00001101100101";
		Trees_din <= x"020f1920";
		wait for Clk_period;
		Addr <=  "00001101100110";
		Trees_din <= x"02030104";
		wait for Clk_period;
		Addr <=  "00001101100111";
		Trees_din <= x"ff960de9";
		wait for Clk_period;
		Addr <=  "00001101101000";
		Trees_din <= x"04ff070c";
		wait for Clk_period;
		Addr <=  "00001101101001";
		Trees_din <= x"08005308";
		wait for Clk_period;
		Addr <=  "00001101101010";
		Trees_din <= x"0bfead04";
		wait for Clk_period;
		Addr <=  "00001101101011";
		Trees_din <= x"005b0de9";
		wait for Clk_period;
		Addr <=  "00001101101100";
		Trees_din <= x"00120de9";
		wait for Clk_period;
		Addr <=  "00001101101101";
		Trees_din <= x"ffe50de9";
		wait for Clk_period;
		Addr <=  "00001101101110";
		Trees_din <= x"08005a0c";
		wait for Clk_period;
		Addr <=  "00001101101111";
		Trees_din <= x"03fbeb04";
		wait for Clk_period;
		Addr <=  "00001101110000";
		Trees_din <= x"00010de9";
		wait for Clk_period;
		Addr <=  "00001101110001";
		Trees_din <= x"06fdbb04";
		wait for Clk_period;
		Addr <=  "00001101110010";
		Trees_din <= x"ffe60de9";
		wait for Clk_period;
		Addr <=  "00001101110011";
		Trees_din <= x"ffa40de9";
		wait for Clk_period;
		Addr <=  "00001101110100";
		Trees_din <= x"001b0de9";
		wait for Clk_period;
		Addr <=  "00001101110101";
		Trees_din <= x"060e1c08";
		wait for Clk_period;
		Addr <=  "00001101110110";
		Trees_din <= x"09fa3b04";
		wait for Clk_period;
		Addr <=  "00001101110111";
		Trees_din <= x"001d0de9";
		wait for Clk_period;
		Addr <=  "00001101111000";
		Trees_din <= x"00690de9";
		wait for Clk_period;
		Addr <=  "00001101111001";
		Trees_din <= x"fff70de9";
		wait for Clk_period;
		Addr <=  "00001101111010";
		Trees_din <= x"02083610";
		wait for Clk_period;
		Addr <=  "00001101111011";
		Trees_din <= x"13028708";
		wait for Clk_period;
		Addr <=  "00001101111100";
		Trees_din <= x"03fbeb04";
		wait for Clk_period;
		Addr <=  "00001101111101";
		Trees_din <= x"ffe70e35";
		wait for Clk_period;
		Addr <=  "00001101111110";
		Trees_din <= x"ff930e35";
		wait for Clk_period;
		Addr <=  "00001101111111";
		Trees_din <= x"08005204";
		wait for Clk_period;
		Addr <=  "00001110000000";
		Trees_din <= x"00320e35";
		wait for Clk_period;
		Addr <=  "00001110000001";
		Trees_din <= x"ffd20e35";
		wait for Clk_period;
		Addr <=  "00001110000010";
		Trees_din <= x"02117810";
		wait for Clk_period;
		Addr <=  "00001110000011";
		Trees_din <= x"04025208";
		wait for Clk_period;
		Addr <=  "00001110000100";
		Trees_din <= x"0c009604";
		wait for Clk_period;
		Addr <=  "00001110000101";
		Trees_din <= x"00020e35";
		wait for Clk_period;
		Addr <=  "00001110000110";
		Trees_din <= x"00410e35";
		wait for Clk_period;
		Addr <=  "00001110000111";
		Trees_din <= x"09027b04";
		wait for Clk_period;
		Addr <=  "00001110001000";
		Trees_din <= x"ffc70e35";
		wait for Clk_period;
		Addr <=  "00001110001001";
		Trees_din <= x"00020e35";
		wait for Clk_period;
		Addr <=  "00001110001010";
		Trees_din <= x"0302e404";
		wait for Clk_period;
		Addr <=  "00001110001011";
		Trees_din <= x"00600e35";
		wait for Clk_period;
		Addr <=  "00001110001100";
		Trees_din <= x"001b0e35";
		wait for Clk_period;
		Addr <=  "00001110001101";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00001110001110";
		Trees_din <= x"020b1e14";
		wait for Clk_period;
		Addr <=  "00001110001111";
		Trees_din <= x"07005908";
		wait for Clk_period;
		Addr <=  "00001110010000";
		Trees_din <= x"04fee804";
		wait for Clk_period;
		Addr <=  "00001110010001";
		Trees_din <= x"ffe60e7d";
		wait for Clk_period;
		Addr <=  "00001110010010";
		Trees_din <= x"ff9c0e7d";
		wait for Clk_period;
		Addr <=  "00001110010011";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00001110010100";
		Trees_din <= x"003d0e7d";
		wait for Clk_period;
		Addr <=  "00001110010101";
		Trees_din <= x"14026704";
		wait for Clk_period;
		Addr <=  "00001110010110";
		Trees_din <= x"ffce0e7d";
		wait for Clk_period;
		Addr <=  "00001110010111";
		Trees_din <= x"fff60e7d";
		wait for Clk_period;
		Addr <=  "00001110011000";
		Trees_din <= x"04081e08";
		wait for Clk_period;
		Addr <=  "00001110011001";
		Trees_din <= x"1b00b704";
		wait for Clk_period;
		Addr <=  "00001110011010";
		Trees_din <= x"00070e7d";
		wait for Clk_period;
		Addr <=  "00001110011011";
		Trees_din <= x"00530e7d";
		wait for Clk_period;
		Addr <=  "00001110011100";
		Trees_din <= x"021ddb04";
		wait for Clk_period;
		Addr <=  "00001110011101";
		Trees_din <= x"ffc30e7d";
		wait for Clk_period;
		Addr <=  "00001110011110";
		Trees_din <= x"00520e7d";
		wait for Clk_period;
		Addr <=  "00001110011111";
		Trees_din <= x"020f1918";
		wait for Clk_period;
		Addr <=  "00001110100000";
		Trees_din <= x"02030104";
		wait for Clk_period;
		Addr <=  "00001110100001";
		Trees_din <= x"ffa40ec1";
		wait for Clk_period;
		Addr <=  "00001110100010";
		Trees_din <= x"01fcdb08";
		wait for Clk_period;
		Addr <=  "00001110100011";
		Trees_din <= x"01fbb404";
		wait for Clk_period;
		Addr <=  "00001110100100";
		Trees_din <= x"fff10ec1";
		wait for Clk_period;
		Addr <=  "00001110100101";
		Trees_din <= x"00470ec1";
		wait for Clk_period;
		Addr <=  "00001110100110";
		Trees_din <= x"18003404";
		wait for Clk_period;
		Addr <=  "00001110100111";
		Trees_din <= x"000d0ec1";
		wait for Clk_period;
		Addr <=  "00001110101000";
		Trees_din <= x"03fb8804";
		wait for Clk_period;
		Addr <=  "00001110101001";
		Trees_din <= x"00070ec1";
		wait for Clk_period;
		Addr <=  "00001110101010";
		Trees_din <= x"ffaf0ec1";
		wait for Clk_period;
		Addr <=  "00001110101011";
		Trees_din <= x"00ce5b08";
		wait for Clk_period;
		Addr <=  "00001110101100";
		Trees_din <= x"021ddb04";
		wait for Clk_period;
		Addr <=  "00001110101101";
		Trees_din <= x"ffdb0ec1";
		wait for Clk_period;
		Addr <=  "00001110101110";
		Trees_din <= x"00500ec1";
		wait for Clk_period;
		Addr <=  "00001110101111";
		Trees_din <= x"00580ec1";
		wait for Clk_period;
		Addr <=  "00001110110000";
		Trees_din <= x"02107418";
		wait for Clk_period;
		Addr <=  "00001110110001";
		Trees_din <= x"0700590c";
		wait for Clk_period;
		Addr <=  "00001110110010";
		Trees_din <= x"020b1e08";
		wait for Clk_period;
		Addr <=  "00001110110011";
		Trees_din <= x"1403b404";
		wait for Clk_period;
		Addr <=  "00001110110100";
		Trees_din <= x"ffaa0efd";
		wait for Clk_period;
		Addr <=  "00001110110101";
		Trees_din <= x"fff00efd";
		wait for Clk_period;
		Addr <=  "00001110110110";
		Trees_din <= x"fff80efd";
		wait for Clk_period;
		Addr <=  "00001110110111";
		Trees_din <= x"17004308";
		wait for Clk_period;
		Addr <=  "00001110111000";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00001110111001";
		Trees_din <= x"00490efd";
		wait for Clk_period;
		Addr <=  "00001110111010";
		Trees_din <= x"00030efd";
		wait for Clk_period;
		Addr <=  "00001110111011";
		Trees_din <= x"ffdc0efd";
		wait for Clk_period;
		Addr <=  "00001110111100";
		Trees_din <= x"0216d904";
		wait for Clk_period;
		Addr <=  "00001110111101";
		Trees_din <= x"00170efd";
		wait for Clk_period;
		Addr <=  "00001110111110";
		Trees_din <= x"00530efd";
		wait for Clk_period;
		Addr <=  "00001110111111";
		Trees_din <= x"020f1918";
		wait for Clk_period;
		Addr <=  "00001111000000";
		Trees_din <= x"0700590c";
		wait for Clk_period;
		Addr <=  "00001111000001";
		Trees_din <= x"04fee804";
		wait for Clk_period;
		Addr <=  "00001111000010";
		Trees_din <= x"fff80f39";
		wait for Clk_period;
		Addr <=  "00001111000011";
		Trees_din <= x"020b1e04";
		wait for Clk_period;
		Addr <=  "00001111000100";
		Trees_din <= x"ffaa0f39";
		wait for Clk_period;
		Addr <=  "00001111000101";
		Trees_din <= x"ffed0f39";
		wait for Clk_period;
		Addr <=  "00001111000110";
		Trees_din <= x"17004308";
		wait for Clk_period;
		Addr <=  "00001111000111";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00001111001000";
		Trees_din <= x"00440f39";
		wait for Clk_period;
		Addr <=  "00001111001001";
		Trees_din <= x"00030f39";
		wait for Clk_period;
		Addr <=  "00001111001010";
		Trees_din <= x"ffd90f39";
		wait for Clk_period;
		Addr <=  "00001111001011";
		Trees_din <= x"00c02704";
		wait for Clk_period;
		Addr <=  "00001111001100";
		Trees_din <= x"00120f39";
		wait for Clk_period;
		Addr <=  "00001111001101";
		Trees_din <= x"004e0f39";
		wait for Clk_period;
		Addr <=  "00001111001110";
		Trees_din <= x"0208360c";
		wait for Clk_period;
		Addr <=  "00001111001111";
		Trees_din <= x"0a000f04";
		wait for Clk_period;
		Addr <=  "00001111010000";
		Trees_din <= x"000f0f7d";
		wait for Clk_period;
		Addr <=  "00001111010001";
		Trees_din <= x"06009f04";
		wait for Clk_period;
		Addr <=  "00001111010010";
		Trees_din <= x"ffa20f7d";
		wait for Clk_period;
		Addr <=  "00001111010011";
		Trees_din <= x"fffa0f7d";
		wait for Clk_period;
		Addr <=  "00001111010100";
		Trees_din <= x"0216d914";
		wait for Clk_period;
		Addr <=  "00001111010101";
		Trees_din <= x"00df9f04";
		wait for Clk_period;
		Addr <=  "00001111010110";
		Trees_din <= x"ffc20f7d";
		wait for Clk_period;
		Addr <=  "00001111010111";
		Trees_din <= x"0a03450c";
		wait for Clk_period;
		Addr <=  "00001111011000";
		Trees_din <= x"020d6208";
		wait for Clk_period;
		Addr <=  "00001111011001";
		Trees_din <= x"16003204";
		wait for Clk_period;
		Addr <=  "00001111011010";
		Trees_din <= x"00270f7d";
		wait for Clk_period;
		Addr <=  "00001111011011";
		Trees_din <= x"ffff0f7d";
		wait for Clk_period;
		Addr <=  "00001111011100";
		Trees_din <= x"004c0f7d";
		wait for Clk_period;
		Addr <=  "00001111011101";
		Trees_din <= x"ffea0f7d";
		wait for Clk_period;
		Addr <=  "00001111011110";
		Trees_din <= x"004d0f7d";
		wait for Clk_period;
		Addr <=  "00001111011111";
		Trees_din <= x"02117818";
		wait for Clk_period;
		Addr <=  "00001111100000";
		Trees_din <= x"03fd9410";
		wait for Clk_period;
		Addr <=  "00001111100001";
		Trees_din <= x"07005808";
		wait for Clk_period;
		Addr <=  "00001111100010";
		Trees_din <= x"09028204";
		wait for Clk_period;
		Addr <=  "00001111100011";
		Trees_din <= x"ffd50fb1";
		wait for Clk_period;
		Addr <=  "00001111100100";
		Trees_din <= x"fffa0fb1";
		wait for Clk_period;
		Addr <=  "00001111100101";
		Trees_din <= x"14018504";
		wait for Clk_period;
		Addr <=  "00001111100110";
		Trees_din <= x"fffc0fb1";
		wait for Clk_period;
		Addr <=  "00001111100111";
		Trees_din <= x"00360fb1";
		wait for Clk_period;
		Addr <=  "00001111101000";
		Trees_din <= x"01fc3604";
		wait for Clk_period;
		Addr <=  "00001111101001";
		Trees_din <= x"fff70fb1";
		wait for Clk_period;
		Addr <=  "00001111101010";
		Trees_din <= x"ffb80fb1";
		wait for Clk_period;
		Addr <=  "00001111101011";
		Trees_din <= x"003f0fb1";
		wait for Clk_period;
		Addr <=  "00001111101100";
		Trees_din <= x"0208360c";
		wait for Clk_period;
		Addr <=  "00001111101101";
		Trees_din <= x"0a000f04";
		wait for Clk_period;
		Addr <=  "00001111101110";
		Trees_din <= x"000d0fed";
		wait for Clk_period;
		Addr <=  "00001111101111";
		Trees_din <= x"03fbf704";
		wait for Clk_period;
		Addr <=  "00001111110000";
		Trees_din <= x"fff00fed";
		wait for Clk_period;
		Addr <=  "00001111110001";
		Trees_din <= x"ffa70fed";
		wait for Clk_period;
		Addr <=  "00001111110010";
		Trees_din <= x"07005a10";
		wait for Clk_period;
		Addr <=  "00001111110011";
		Trees_din <= x"020fd908";
		wait for Clk_period;
		Addr <=  "00001111110100";
		Trees_din <= x"10011f04";
		wait for Clk_period;
		Addr <=  "00001111110101";
		Trees_din <= x"ffd30fed";
		wait for Clk_period;
		Addr <=  "00001111110110";
		Trees_din <= x"000a0fed";
		wait for Clk_period;
		Addr <=  "00001111110111";
		Trees_din <= x"03015d04";
		wait for Clk_period;
		Addr <=  "00001111111000";
		Trees_din <= x"00390fed";
		wait for Clk_period;
		Addr <=  "00001111111001";
		Trees_din <= x"00030fed";
		wait for Clk_period;
		Addr <=  "00001111111010";
		Trees_din <= x"00430fed";
		wait for Clk_period;
		Addr <=  "00001111111011";
		Trees_din <= x"02083608";
		wait for Clk_period;
		Addr <=  "00001111111100";
		Trees_din <= x"13028704";
		wait for Clk_period;
		Addr <=  "00001111111101";
		Trees_din <= x"ffb91021";
		wait for Clk_period;
		Addr <=  "00001111111110";
		Trees_din <= x"00071021";
		wait for Clk_period;
		Addr <=  "00001111111111";
		Trees_din <= x"0216d910";
		wait for Clk_period;
		Addr <=  "00010000000000";
		Trees_din <= x"00eab204";
		wait for Clk_period;
		Addr <=  "00010000000001";
		Trees_din <= x"ffd31021";
		wait for Clk_period;
		Addr <=  "00010000000010";
		Trees_din <= x"0fff2e04";
		wait for Clk_period;
		Addr <=  "00010000000011";
		Trees_din <= x"fff41021";
		wait for Clk_period;
		Addr <=  "00010000000100";
		Trees_din <= x"11029104";
		wait for Clk_period;
		Addr <=  "00010000000101";
		Trees_din <= x"003b1021";
		wait for Clk_period;
		Addr <=  "00010000000110";
		Trees_din <= x"00101021";
		wait for Clk_period;
		Addr <=  "00010000000111";
		Trees_din <= x"00431021";
		wait for Clk_period;
		Addr <=  "00010000001000";
		Trees_din <= x"020f1910";
		wait for Clk_period;
		Addr <=  "00010000001001";
		Trees_din <= x"1700440c";
		wait for Clk_period;
		Addr <=  "00010000001010";
		Trees_din <= x"17004208";
		wait for Clk_period;
		Addr <=  "00010000001011";
		Trees_din <= x"18003404";
		wait for Clk_period;
		Addr <=  "00010000001100";
		Trees_din <= x"0001104d";
		wait for Clk_period;
		Addr <=  "00010000001101";
		Trees_din <= x"ffcf104d";
		wait for Clk_period;
		Addr <=  "00010000001110";
		Trees_din <= x"0033104d";
		wait for Clk_period;
		Addr <=  "00010000001111";
		Trees_din <= x"ffc9104d";
		wait for Clk_period;
		Addr <=  "00010000010000";
		Trees_din <= x"00c02704";
		wait for Clk_period;
		Addr <=  "00010000010001";
		Trees_din <= x"000c104d";
		wait for Clk_period;
		Addr <=  "00010000010010";
		Trees_din <= x"0041104d";
		wait for Clk_period;
		Addr <=  "00010000010011";
		Trees_din <= x"02083608";
		wait for Clk_period;
		Addr <=  "00010000010100";
		Trees_din <= x"13028704";
		wait for Clk_period;
		Addr <=  "00010000010101";
		Trees_din <= x"ffbf1079";
		wait for Clk_period;
		Addr <=  "00010000010110";
		Trees_din <= x"00041079";
		wait for Clk_period;
		Addr <=  "00010000010111";
		Trees_din <= x"07005a0c";
		wait for Clk_period;
		Addr <=  "00010000011000";
		Trees_din <= x"02159b08";
		wait for Clk_period;
		Addr <=  "00010000011001";
		Trees_din <= x"04025204";
		wait for Clk_period;
		Addr <=  "00010000011010";
		Trees_din <= x"000e1079";
		wait for Clk_period;
		Addr <=  "00010000011011";
		Trees_din <= x"ffd31079";
		wait for Clk_period;
		Addr <=  "00010000011100";
		Trees_din <= x"002b1079";
		wait for Clk_period;
		Addr <=  "00010000011101";
		Trees_din <= x"003d1079";
		wait for Clk_period;
		Addr <=  "00010000011110";
		Trees_din <= x"020b1e10";
		wait for Clk_period;
		Addr <=  "00010000011111";
		Trees_din <= x"07005908";
		wait for Clk_period;
		Addr <=  "00010000100000";
		Trees_din <= x"04fee804";
		wait for Clk_period;
		Addr <=  "00010000100001";
		Trees_din <= x"fff110ad";
		wait for Clk_period;
		Addr <=  "00010000100010";
		Trees_din <= x"ffb710ad";
		wait for Clk_period;
		Addr <=  "00010000100011";
		Trees_din <= x"07005a04";
		wait for Clk_period;
		Addr <=  "00010000100100";
		Trees_din <= x"002110ad";
		wait for Clk_period;
		Addr <=  "00010000100101";
		Trees_din <= x"ffe410ad";
		wait for Clk_period;
		Addr <=  "00010000100110";
		Trees_din <= x"0fff2e04";
		wait for Clk_period;
		Addr <=  "00010000100111";
		Trees_din <= x"fff710ad";
		wait for Clk_period;
		Addr <=  "00010000101000";
		Trees_din <= x"09fb1604";
		wait for Clk_period;
		Addr <=  "00010000101001";
		Trees_din <= x"000110ad";
		wait for Clk_period;
		Addr <=  "00010000101010";
		Trees_din <= x"004410ad";
		wait for Clk_period;
		Addr <=  "00010000101011";
		Trees_din <= x"02117810";
		wait for Clk_period;
		Addr <=  "00010000101100";
		Trees_din <= x"0400750c";
		wait for Clk_period;
		Addr <=  "00010000101101";
		Trees_din <= x"05058708";
		wait for Clk_period;
		Addr <=  "00010000101110";
		Trees_din <= x"15028704";
		wait for Clk_period;
		Addr <=  "00010000101111";
		Trees_din <= x"fffb10d1";
		wait for Clk_period;
		Addr <=  "00010000110000";
		Trees_din <= x"003010d1";
		wait for Clk_period;
		Addr <=  "00010000110001";
		Trees_din <= x"ffde10d1";
		wait for Clk_period;
		Addr <=  "00010000110010";
		Trees_din <= x"ffcf10d1";
		wait for Clk_period;
		Addr <=  "00010000110011";
		Trees_din <= x"003110d1";
		wait for Clk_period;
		Addr <=  "00010000110100";
		Trees_din <= x"020b1e08";
		wait for Clk_period;
		Addr <=  "00010000110101";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00010000110110";
		Trees_din <= x"ffc910f5";
		wait for Clk_period;
		Addr <=  "00010000110111";
		Trees_din <= x"000210f5";
		wait for Clk_period;
		Addr <=  "00010000111000";
		Trees_din <= x"04081e08";
		wait for Clk_period;
		Addr <=  "00010000111001";
		Trees_din <= x"1b017204";
		wait for Clk_period;
		Addr <=  "00010000111010";
		Trees_din <= x"000510f5";
		wait for Clk_period;
		Addr <=  "00010000111011";
		Trees_din <= x"004210f5";
		wait for Clk_period;
		Addr <=  "00010000111100";
		Trees_din <= x"fffb10f5";
		wait for Clk_period;
		Addr <=  "00010000111101";
		Trees_din <= x"0216d914";
		wait for Clk_period;
		Addr <=  "00010000111110";
		Trees_din <= x"03fd940c";
		wait for Clk_period;
		Addr <=  "00010000111111";
		Trees_din <= x"02069704";
		wait for Clk_period;
		Addr <=  "00010001000000";
		Trees_din <= x"ffe51121";
		wait for Clk_period;
		Addr <=  "00010001000001";
		Trees_din <= x"18003a04";
		wait for Clk_period;
		Addr <=  "00010001000010";
		Trees_din <= x"fffd1121";
		wait for Clk_period;
		Addr <=  "00010001000011";
		Trees_din <= x"00341121";
		wait for Clk_period;
		Addr <=  "00010001000100";
		Trees_din <= x"13027a04";
		wait for Clk_period;
		Addr <=  "00010001000101";
		Trees_din <= x"ffc41121";
		wait for Clk_period;
		Addr <=  "00010001000110";
		Trees_din <= x"fff81121";
		wait for Clk_period;
		Addr <=  "00010001000111";
		Trees_din <= x"00391121";
		wait for Clk_period;
		Addr <=  "00010001001000";
		Trees_din <= x"020b1e0c";
		wait for Clk_period;
		Addr <=  "00010001001001";
		Trees_din <= x"0a001604";
		wait for Clk_period;
		Addr <=  "00010001001010";
		Trees_din <= x"000a114d";
		wait for Clk_period;
		Addr <=  "00010001001011";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00010001001100";
		Trees_din <= x"ffc0114d";
		wait for Clk_period;
		Addr <=  "00010001001101";
		Trees_din <= x"fff7114d";
		wait for Clk_period;
		Addr <=  "00010001001110";
		Trees_din <= x"0fff2e04";
		wait for Clk_period;
		Addr <=  "00010001001111";
		Trees_din <= x"fff7114d";
		wait for Clk_period;
		Addr <=  "00010001010000";
		Trees_din <= x"09fb1604";
		wait for Clk_period;
		Addr <=  "00010001010001";
		Trees_din <= x"ffff114d";
		wait for Clk_period;
		Addr <=  "00010001010010";
		Trees_din <= x"003e114d";
		wait for Clk_period;
		Addr <=  "00010001010011";
		Trees_din <= x"02159b10";
		wait for Clk_period;
		Addr <=  "00010001010100";
		Trees_din <= x"03fd9408";
		wait for Clk_period;
		Addr <=  "00010001010101";
		Trees_din <= x"18003904";
		wait for Clk_period;
		Addr <=  "00010001010110";
		Trees_din <= x"ffef1171";
		wait for Clk_period;
		Addr <=  "00010001010111";
		Trees_din <= x"001e1171";
		wait for Clk_period;
		Addr <=  "00010001011000";
		Trees_din <= x"12009804";
		wait for Clk_period;
		Addr <=  "00010001011001";
		Trees_din <= x"ffbf1171";
		wait for Clk_period;
		Addr <=  "00010001011010";
		Trees_din <= x"fff71171";
		wait for Clk_period;
		Addr <=  "00010001011011";
		Trees_din <= x"00331171";
		wait for Clk_period;
		Addr <=  "00010001011100";
		Trees_din <= x"02088f08";
		wait for Clk_period;
		Addr <=  "00010001011101";
		Trees_din <= x"01fcd504";
		wait for Clk_period;
		Addr <=  "00010001011110";
		Trees_din <= x"00001195";
		wait for Clk_period;
		Addr <=  "00010001011111";
		Trees_din <= x"ffc71195";
		wait for Clk_period;
		Addr <=  "00010001100000";
		Trees_din <= x"07005a08";
		wait for Clk_period;
		Addr <=  "00010001100001";
		Trees_din <= x"0c00dd04";
		wait for Clk_period;
		Addr <=  "00010001100010";
		Trees_din <= x"ffea1195";
		wait for Clk_period;
		Addr <=  "00010001100011";
		Trees_din <= x"001a1195";
		wait for Clk_period;
		Addr <=  "00010001100100";
		Trees_din <= x"00341195";
		wait for Clk_period;
		Addr <=  "00010001100101";
		Trees_din <= x"020b1e0c";
		wait for Clk_period;
		Addr <=  "00010001100110";
		Trees_din <= x"0a001604";
		wait for Clk_period;
		Addr <=  "00010001100111";
		Trees_din <= x"000911c1";
		wait for Clk_period;
		Addr <=  "00010001101000";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00010001101001";
		Trees_din <= x"ffc511c1";
		wait for Clk_period;
		Addr <=  "00010001101010";
		Trees_din <= x"fff611c1";
		wait for Clk_period;
		Addr <=  "00010001101011";
		Trees_din <= x"10fffc04";
		wait for Clk_period;
		Addr <=  "00010001101100";
		Trees_din <= x"fffa11c1";
		wait for Clk_period;
		Addr <=  "00010001101101";
		Trees_din <= x"09feb404";
		wait for Clk_period;
		Addr <=  "00010001101110";
		Trees_din <= x"000f11c1";
		wait for Clk_period;
		Addr <=  "00010001101111";
		Trees_din <= x"003511c1";
		wait for Clk_period;
		Addr <=  "00010001110000";
		Trees_din <= x"02088f08";
		wait for Clk_period;
		Addr <=  "00010001110001";
		Trees_din <= x"01fcd504";
		wait for Clk_period;
		Addr <=  "00010001110010";
		Trees_din <= x"000011e5";
		wait for Clk_period;
		Addr <=  "00010001110011";
		Trees_din <= x"ffcc11e5";
		wait for Clk_period;
		Addr <=  "00010001110100";
		Trees_din <= x"0a032a08";
		wait for Clk_period;
		Addr <=  "00010001110101";
		Trees_din <= x"04081e04";
		wait for Clk_period;
		Addr <=  "00010001110110";
		Trees_din <= x"002e11e5";
		wait for Clk_period;
		Addr <=  "00010001110111";
		Trees_din <= x"ffff11e5";
		wait for Clk_period;
		Addr <=  "00010001111000";
		Trees_din <= x"fff211e5";
		wait for Clk_period;
		Addr <=  "00010001111001";
		Trees_din <= x"020b1e08";
		wait for Clk_period;
		Addr <=  "00010001111010";
		Trees_din <= x"00097504";
		wait for Clk_period;
		Addr <=  "00010001111011";
		Trees_din <= x"ffd21201";
		wait for Clk_period;
		Addr <=  "00010001111100";
		Trees_din <= x"00061201";
		wait for Clk_period;
		Addr <=  "00010001111101";
		Trees_din <= x"10fffc04";
		wait for Clk_period;
		Addr <=  "00010001111110";
		Trees_din <= x"fffa1201";
		wait for Clk_period;
		Addr <=  "00010001111111";
		Trees_din <= x"00271201";
		wait for Clk_period;
		Addr <=  "00010010000000";
		Trees_din <= x"0216d910";
		wait for Clk_period;
		Addr <=  "00010010000001";
		Trees_din <= x"03fd9408";
		wait for Clk_period;
		Addr <=  "00010010000010";
		Trees_din <= x"07005804";
		wait for Clk_period;
		Addr <=  "00010010000011";
		Trees_din <= x"fff11225";
		wait for Clk_period;
		Addr <=  "00010010000100";
		Trees_din <= x"001c1225";
		wait for Clk_period;
		Addr <=  "00010010000101";
		Trees_din <= x"13021e04";
		wait for Clk_period;
		Addr <=  "00010010000110";
		Trees_din <= x"ffca1225";
		wait for Clk_period;
		Addr <=  "00010010000111";
		Trees_din <= x"fff41225";
		wait for Clk_period;
		Addr <=  "00010010001000";
		Trees_din <= x"00311225";
		wait for Clk_period;
		Addr <=  "00010010001001";
		Trees_din <= x"02056d04";
		wait for Clk_period;
		Addr <=  "00010010001010";
		Trees_din <= x"ffd71241";
		wait for Clk_period;
		Addr <=  "00010010001011";
		Trees_din <= x"0a032a08";
		wait for Clk_period;
		Addr <=  "00010010001100";
		Trees_din <= x"16007d04";
		wait for Clk_period;
		Addr <=  "00010010001101";
		Trees_din <= x"002d1241";
		wait for Clk_period;
		Addr <=  "00010010001110";
		Trees_din <= x"00001241";
		wait for Clk_period;
		Addr <=  "00010010001111";
		Trees_din <= x"ffee1241";
		wait for Clk_period;
		Addr <=  "00010010010000";
		Trees_din <= x"020b1e08";
		wait for Clk_period;
		Addr <=  "00010010010001";
		Trees_din <= x"03fbf704";
		wait for Clk_period;
		Addr <=  "00010010010010";
		Trees_din <= x"00071265";
		wait for Clk_period;
		Addr <=  "00010010010011";
		Trees_din <= x"ffd51265";
		wait for Clk_period;
		Addr <=  "00010010010100";
		Trees_din <= x"04081e08";
		wait for Clk_period;
		Addr <=  "00010010010101";
		Trees_din <= x"15043104";
		wait for Clk_period;
		Addr <=  "00010010010110";
		Trees_din <= x"00341265";
		wait for Clk_period;
		Addr <=  "00010010010111";
		Trees_din <= x"00041265";
		wait for Clk_period;
		Addr <=  "00010010011000";
		Trees_din <= x"fff91265";
		wait for Clk_period;
		Addr <=  "00010010011001";
		Trees_din <= x"02056d04";
		wait for Clk_period;
		Addr <=  "00010010011010";
		Trees_din <= x"ffdc1289";
		wait for Clk_period;
		Addr <=  "00010010011011";
		Trees_din <= x"0a032a0c";
		wait for Clk_period;
		Addr <=  "00010010011100";
		Trees_din <= x"11031a08";
		wait for Clk_period;
		Addr <=  "00010010011101";
		Trees_din <= x"03fe3304";
		wait for Clk_period;
		Addr <=  "00010010011110";
		Trees_din <= x"002f1289";
		wait for Clk_period;
		Addr <=  "00010010011111";
		Trees_din <= x"00081289";
		wait for Clk_period;
		Addr <=  "00010010100000";
		Trees_din <= x"fffa1289";
		wait for Clk_period;
		Addr <=  "00010010100001";
		Trees_din <= x"ffef1289";
		wait for Clk_period;
		Addr <=  "00010010100010";
		Trees_din <= x"020b1e08";
		wait for Clk_period;
		Addr <=  "00010010100011";
		Trees_din <= x"00097504";
		wait for Clk_period;
		Addr <=  "00010010100100";
		Trees_din <= x"ffd612a5";
		wait for Clk_period;
		Addr <=  "00010010100101";
		Trees_din <= x"000912a5";
		wait for Clk_period;
		Addr <=  "00010010100110";
		Trees_din <= x"09fdbe04";
		wait for Clk_period;
		Addr <=  "00010010100111";
		Trees_din <= x"fffb12a5";
		wait for Clk_period;
		Addr <=  "00010010101000";
		Trees_din <= x"002512a5";
		wait for Clk_period;
		Addr <=  "00010010101001";
		Trees_din <= x"02056d04";
		wait for Clk_period;
		Addr <=  "00010010101010";
		Trees_din <= x"ffdf12c1";
		wait for Clk_period;
		Addr <=  "00010010101011";
		Trees_din <= x"0a032a08";
		wait for Clk_period;
		Addr <=  "00010010101100";
		Trees_din <= x"16007d04";
		wait for Clk_period;
		Addr <=  "00010010101101";
		Trees_din <= x"002712c1";
		wait for Clk_period;
		Addr <=  "00010010101110";
		Trees_din <= x"000012c1";
		wait for Clk_period;
		Addr <=  "00010010101111";
		Trees_din <= x"fff112c1";
		wait for Clk_period;
		Addr <=  "00010010110000";
		Trees_din <= x"020b1e08";
		wait for Clk_period;
		Addr <=  "00010010110001";
		Trees_din <= x"03fbf704";
		wait for Clk_period;
		Addr <=  "00010010110010";
		Trees_din <= x"000a12dd";
		wait for Clk_period;
		Addr <=  "00010010110011";
		Trees_din <= x"ffd912dd";
		wait for Clk_period;
		Addr <=  "00010010110100";
		Trees_din <= x"10fffc04";
		wait for Clk_period;
		Addr <=  "00010010110101";
		Trees_din <= x"fff712dd";
		wait for Clk_period;
		Addr <=  "00010010110110";
		Trees_din <= x"002012dd";
		wait for Clk_period;
		Addr <=  "00010010110111";
		Trees_din <= x"02056d04";
		wait for Clk_period;
		Addr <=  "00010010111000";
		Trees_din <= x"ffe21301";
		wait for Clk_period;
		Addr <=  "00010010111001";
		Trees_din <= x"03fdb908";
		wait for Clk_period;
		Addr <=  "00010010111010";
		Trees_din <= x"1c003504";
		wait for Clk_period;
		Addr <=  "00010010111011";
		Trees_din <= x"00281301";
		wait for Clk_period;
		Addr <=  "00010010111100";
		Trees_din <= x"00041301";
		wait for Clk_period;
		Addr <=  "00010010111101";
		Trees_din <= x"16002c04";
		wait for Clk_period;
		Addr <=  "00010010111110";
		Trees_din <= x"000b1301";
		wait for Clk_period;
		Addr <=  "00010010111111";
		Trees_din <= x"ffe91301";
		wait for Clk_period;
		Addr <=  "00010011000000";
		Trees_din <= x"020b1e08";
		wait for Clk_period;
		Addr <=  "00010011000001";
		Trees_din <= x"00097504";
		wait for Clk_period;
		Addr <=  "00010011000010";
		Trees_din <= x"ffda131d";
		wait for Clk_period;
		Addr <=  "00010011000011";
		Trees_din <= x"000a131d";
		wait for Clk_period;
		Addr <=  "00010011000100";
		Trees_din <= x"04081e04";
		wait for Clk_period;
		Addr <=  "00010011000101";
		Trees_din <= x"001f131d";
		wait for Clk_period;
		Addr <=  "00010011000110";
		Trees_din <= x"fff8131d";
		wait for Clk_period;
		Addr <=  "00010011000111";
		Trees_din <= x"1700440c";
		wait for Clk_period;
		Addr <=  "00010011001000";
		Trees_din <= x"1c003004";
		wait for Clk_period;
		Addr <=  "00010011001001";
		Trees_din <= x"ffe61341";
		wait for Clk_period;
		Addr <=  "00010011001010";
		Trees_din <= x"0c015304";
		wait for Clk_period;
		Addr <=  "00010011001011";
		Trees_din <= x"000e1341";
		wait for Clk_period;
		Addr <=  "00010011001100";
		Trees_din <= x"00301341";
		wait for Clk_period;
		Addr <=  "00010011001101";
		Trees_din <= x"09028804";
		wait for Clk_period;
		Addr <=  "00010011001110";
		Trees_din <= x"ffdc1341";
		wait for Clk_period;
		Addr <=  "00010011001111";
		Trees_din <= x"00021341";
		wait for Clk_period;
		Addr <=  "00010011010000";
		Trees_din <= x"020b1e08";
		wait for Clk_period;
		Addr <=  "00010011010001";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00010011010010";
		Trees_din <= x"ffd9135d";
		wait for Clk_period;
		Addr <=  "00010011010011";
		Trees_din <= x"0009135d";
		wait for Clk_period;
		Addr <=  "00010011010100";
		Trees_din <= x"10fffc04";
		wait for Clk_period;
		Addr <=  "00010011010101";
		Trees_din <= x"fff8135d";
		wait for Clk_period;
		Addr <=  "00010011010110";
		Trees_din <= x"001e135d";
		wait for Clk_period;
		Addr <=  "00010011010111";
		Trees_din <= x"02056d04";
		wait for Clk_period;
		Addr <=  "00010011011000";
		Trees_din <= x"ffe31379";
		wait for Clk_period;
		Addr <=  "00010011011001";
		Trees_din <= x"0a032a08";
		wait for Clk_period;
		Addr <=  "00010011011010";
		Trees_din <= x"03fe3304";
		wait for Clk_period;
		Addr <=  "00010011011011";
		Trees_din <= x"00221379";
		wait for Clk_period;
		Addr <=  "00010011011100";
		Trees_din <= x"fffe1379";
		wait for Clk_period;
		Addr <=  "00010011011101";
		Trees_din <= x"fff11379";
		wait for Clk_period;
		Addr <=  "00010011011110";
		Trees_din <= x"020b1e08";
		wait for Clk_period;
		Addr <=  "00010011011111";
		Trees_din <= x"00097504";
		wait for Clk_period;
		Addr <=  "00010011100000";
		Trees_din <= x"ffdc1395";
		wait for Clk_period;
		Addr <=  "00010011100001";
		Trees_din <= x"00091395";
		wait for Clk_period;
		Addr <=  "00010011100010";
		Trees_din <= x"09fdbe04";
		wait for Clk_period;
		Addr <=  "00010011100011";
		Trees_din <= x"fff91395";
		wait for Clk_period;
		Addr <=  "00010011100100";
		Trees_din <= x"001f1395";
		wait for Clk_period;
		Addr <=  "00010011100101";
		Trees_din <= x"17004408";
		wait for Clk_period;
		Addr <=  "00010011100110";
		Trees_din <= x"1c003004";
		wait for Clk_period;
		Addr <=  "00010011100111";
		Trees_din <= x"ffe813a9";
		wait for Clk_period;
		Addr <=  "00010011101000";
		Trees_din <= x"002513a9";
		wait for Clk_period;
		Addr <=  "00010011101001";
		Trees_din <= x"ffeb13a9";
		wait for Clk_period;
		Addr <=  "00010011101010";
		Trees_din <= x"02056d04";
		wait for Clk_period;
		Addr <=  "00010011101011";
		Trees_din <= x"ffe313c5";
		wait for Clk_period;
		Addr <=  "00010011101100";
		Trees_din <= x"0f022208";
		wait for Clk_period;
		Addr <=  "00010011101101";
		Trees_din <= x"18003a04";
		wait for Clk_period;
		Addr <=  "00010011101110";
		Trees_din <= x"ffe913c5";
		wait for Clk_period;
		Addr <=  "00010011101111";
		Trees_din <= x"001013c5";
		wait for Clk_period;
		Addr <=  "00010011110000";
		Trees_din <= x"001913c5";
		wait for Clk_period;
		Addr <=  "00010011110001";
		Trees_din <= x"020b1e08";
		wait for Clk_period;
		Addr <=  "00010011110010";
		Trees_din <= x"03fbf704";
		wait for Clk_period;
		Addr <=  "00010011110011";
		Trees_din <= x"000813e1";
		wait for Clk_period;
		Addr <=  "00010011110100";
		Trees_din <= x"ffde13e1";
		wait for Clk_period;
		Addr <=  "00010011110101";
		Trees_din <= x"09fdbe04";
		wait for Clk_period;
		Addr <=  "00010011110110";
		Trees_din <= x"fffb13e1";
		wait for Clk_period;
		Addr <=  "00010011110111";
		Trees_din <= x"001d13e1";
		wait for Clk_period;
		Addr <=  "00010011111000";
		Trees_din <= x"02083604";
		wait for Clk_period;
		Addr <=  "00010011111001";
		Trees_din <= x"ffeb13f5";
		wait for Clk_period;
		Addr <=  "00010011111010";
		Trees_din <= x"0f01f304";
		wait for Clk_period;
		Addr <=  "00010011111011";
		Trees_din <= x"fff913f5";
		wait for Clk_period;
		Addr <=  "00010011111100";
		Trees_din <= x"001d13f5";
		wait for Clk_period;
		Addr <=  "00010011111101";
		Trees_din <= x"17004408";
		wait for Clk_period;
		Addr <=  "00010011111110";
		Trees_din <= x"1c003004";
		wait for Clk_period;
		Addr <=  "00010011111111";
		Trees_din <= x"ffec1409";
		wait for Clk_period;
		Addr <=  "00010100000000";
		Trees_din <= x"00221409";
		wait for Clk_period;
		Addr <=  "00010100000001";
		Trees_din <= x"ffed1409";
		wait for Clk_period;
		Addr <=  "00010100000010";
		Trees_din <= x"08005408";
		wait for Clk_period;
		Addr <=  "00010100000011";
		Trees_din <= x"04ff8e04";
		wait for Clk_period;
		Addr <=  "00010100000100";
		Trees_din <= x"001f1425";
		wait for Clk_period;
		Addr <=  "00010100000101";
		Trees_din <= x"fffd1425";
		wait for Clk_period;
		Addr <=  "00010100000110";
		Trees_din <= x"08005704";
		wait for Clk_period;
		Addr <=  "00010100000111";
		Trees_din <= x"ffdf1425";
		wait for Clk_period;
		Addr <=  "00010100001000";
		Trees_din <= x"00061425";
		wait for Clk_period;
		Addr <=  "00010100001001";
		Trees_din <= x"020b1e08";
		wait for Clk_period;
		Addr <=  "00010100001010";
		Trees_din <= x"01fcd504";
		wait for Clk_period;
		Addr <=  "00010100001011";
		Trees_din <= x"00081441";
		wait for Clk_period;
		Addr <=  "00010100001100";
		Trees_din <= x"ffde1441";
		wait for Clk_period;
		Addr <=  "00010100001101";
		Trees_din <= x"10fffc04";
		wait for Clk_period;
		Addr <=  "00010100001110";
		Trees_din <= x"fff81441";
		wait for Clk_period;
		Addr <=  "00010100001111";
		Trees_din <= x"001b1441";
		wait for Clk_period;
		Addr <=  "00010100010000";
		Trees_din <= x"09028708";
		wait for Clk_period;
		Addr <=  "00010100010001";
		Trees_din <= x"12009404";
		wait for Clk_period;
		Addr <=  "00010100010010";
		Trees_din <= x"ffe5145d";
		wait for Clk_period;
		Addr <=  "00010100010011";
		Trees_din <= x"0000145d";
		wait for Clk_period;
		Addr <=  "00010100010100";
		Trees_din <= x"0904c904";
		wait for Clk_period;
		Addr <=  "00010100010101";
		Trees_din <= x"001e145d";
		wait for Clk_period;
		Addr <=  "00010100010110";
		Trees_din <= x"fff6145d";
		wait for Clk_period;
		Addr <=  "00010100010111";
		Trees_din <= x"17004408";
		wait for Clk_period;
		Addr <=  "00010100011000";
		Trees_din <= x"1c003004";
		wait for Clk_period;
		Addr <=  "00010100011001";
		Trees_din <= x"ffee1471";
		wait for Clk_period;
		Addr <=  "00010100011010";
		Trees_din <= x"001e1471";
		wait for Clk_period;
		Addr <=  "00010100011011";
		Trees_din <= x"ffef1471";
		wait for Clk_period;
		Addr <=  "00010100011100";
		Trees_din <= x"02069704";
		wait for Clk_period;
		Addr <=  "00010100011101";
		Trees_din <= x"ffe61485";
		wait for Clk_period;
		Addr <=  "00010100011110";
		Trees_din <= x"04025204";
		wait for Clk_period;
		Addr <=  "00010100011111";
		Trees_din <= x"001a1485";
		wait for Clk_period;
		Addr <=  "00010100100000";
		Trees_din <= x"fffb1485";
		wait for Clk_period;
		Addr <=  "00010100100001";
		Trees_din <= x"020b1e08";
		wait for Clk_period;
		Addr <=  "00010100100010";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00010100100011";
		Trees_din <= x"ffde14a1";
		wait for Clk_period;
		Addr <=  "00010100100100";
		Trees_din <= x"000614a1";
		wait for Clk_period;
		Addr <=  "00010100100101";
		Trees_din <= x"08005604";
		wait for Clk_period;
		Addr <=  "00010100100110";
		Trees_din <= x"001c14a1";
		wait for Clk_period;
		Addr <=  "00010100100111";
		Trees_din <= x"fffb14a1";
		wait for Clk_period;
		Addr <=  "00010100101000";
		Trees_din <= x"09028708";
		wait for Clk_period;
		Addr <=  "00010100101001";
		Trees_din <= x"06ffa104";
		wait for Clk_period;
		Addr <=  "00010100101010";
		Trees_din <= x"000014bd";
		wait for Clk_period;
		Addr <=  "00010100101011";
		Trees_din <= x"ffe914bd";
		wait for Clk_period;
		Addr <=  "00010100101100";
		Trees_din <= x"0904c904";
		wait for Clk_period;
		Addr <=  "00010100101101";
		Trees_din <= x"001b14bd";
		wait for Clk_period;
		Addr <=  "00010100101110";
		Trees_din <= x"fff714bd";
		wait for Clk_period;
		Addr <=  "00010100101111";
		Trees_din <= x"08005404";
		wait for Clk_period;
		Addr <=  "00010100110000";
		Trees_din <= x"000f14d1";
		wait for Clk_period;
		Addr <=  "00010100110001";
		Trees_din <= x"08005704";
		wait for Clk_period;
		Addr <=  "00010100110010";
		Trees_din <= x"ffe314d1";
		wait for Clk_period;
		Addr <=  "00010100110011";
		Trees_din <= x"000614d1";
		wait for Clk_period;
		Addr <=  "00010100110100";
		Trees_din <= x"020b1e08";
		wait for Clk_period;
		Addr <=  "00010100110101";
		Trees_din <= x"01fcd504";
		wait for Clk_period;
		Addr <=  "00010100110110";
		Trees_din <= x"000614ed";
		wait for Clk_period;
		Addr <=  "00010100110111";
		Trees_din <= x"ffdf14ed";
		wait for Clk_period;
		Addr <=  "00010100111000";
		Trees_din <= x"15043804";
		wait for Clk_period;
		Addr <=  "00010100111001";
		Trees_din <= x"001b14ed";
		wait for Clk_period;
		Addr <=  "00010100111010";
		Trees_din <= x"fffb14ed";
		wait for Clk_period;
		Addr <=  "00010100111011";
		Trees_din <= x"12009404";
		wait for Clk_period;
		Addr <=  "00010100111100";
		Trees_din <= x"fff01501";
		wait for Clk_period;
		Addr <=  "00010100111101";
		Trees_din <= x"1c003004";
		wait for Clk_period;
		Addr <=  "00010100111110";
		Trees_din <= x"fff31501";
		wait for Clk_period;
		Addr <=  "00010100111111";
		Trees_din <= x"001b1501";
		wait for Clk_period;
		Addr <=  "00010101000000";
		Trees_din <= x"1402cd08";
		wait for Clk_period;
		Addr <=  "00010101000001";
		Trees_din <= x"18003904";
		wait for Clk_period;
		Addr <=  "00010101000010";
		Trees_din <= x"ffe2151d";
		wait for Clk_period;
		Addr <=  "00010101000011";
		Trees_din <= x"000b151d";
		wait for Clk_period;
		Addr <=  "00010101000100";
		Trees_din <= x"1300c004";
		wait for Clk_period;
		Addr <=  "00010101000101";
		Trees_din <= x"ffff151d";
		wait for Clk_period;
		Addr <=  "00010101000110";
		Trees_din <= x"0017151d";
		wait for Clk_period;
		Addr <=  "00010101000111";
		Trees_din <= x"02072404";
		wait for Clk_period;
		Addr <=  "00010101001000";
		Trees_din <= x"ffe71531";
		wait for Clk_period;
		Addr <=  "00010101001001";
		Trees_din <= x"04025204";
		wait for Clk_period;
		Addr <=  "00010101001010";
		Trees_din <= x"001a1531";
		wait for Clk_period;
		Addr <=  "00010101001011";
		Trees_din <= x"fffd1531";
		wait for Clk_period;
		Addr <=  "00010101001100";
		Trees_din <= x"020b1e08";
		wait for Clk_period;
		Addr <=  "00010101001101";
		Trees_din <= x"06fe6a04";
		wait for Clk_period;
		Addr <=  "00010101001110";
		Trees_din <= x"ffe4154d";
		wait for Clk_period;
		Addr <=  "00010101001111";
		Trees_din <= x"0002154d";
		wait for Clk_period;
		Addr <=  "00010101010000";
		Trees_din <= x"04081e04";
		wait for Clk_period;
		Addr <=  "00010101010001";
		Trees_din <= x"001a154d";
		wait for Clk_period;
		Addr <=  "00010101010010";
		Trees_din <= x"fffb154d";
		wait for Clk_period;
		Addr <=  "00010101010011";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  5
        -----------
		Addr <=  "00000000000000";
		Trees_din <= x"040ebb38";
		wait for Clk_period;
		Addr <=  "00000000000001";
		Trees_din <= x"0406af14";
		wait for Clk_period;
		Addr <=  "00000000000010";
		Trees_din <= x"04048f04";
		wait for Clk_period;
		Addr <=  "00000000000011";
		Trees_din <= x"ff4d0095";
		wait for Clk_period;
		Addr <=  "00000000000100";
		Trees_din <= x"00f7bd04";
		wait for Clk_period;
		Addr <=  "00000000000101";
		Trees_din <= x"ff500095";
		wait for Clk_period;
		Addr <=  "00000000000110";
		Trees_din <= x"05fe0a08";
		wait for Clk_period;
		Addr <=  "00000000000111";
		Trees_din <= x"15053604";
		wait for Clk_period;
		Addr <=  "00000000001000";
		Trees_din <= x"ff6c0095";
		wait for Clk_period;
		Addr <=  "00000000001001";
		Trees_din <= x"00270095";
		wait for Clk_period;
		Addr <=  "00000000001010";
		Trees_din <= x"01870095";
		wait for Clk_period;
		Addr <=  "00000000001011";
		Trees_din <= x"00f01314";
		wait for Clk_period;
		Addr <=  "00000000001100";
		Trees_din <= x"00dc8808";
		wait for Clk_period;
		Addr <=  "00000000001101";
		Trees_din <= x"15f73a04";
		wait for Clk_period;
		Addr <=  "00000000001110";
		Trees_din <= x"00120095";
		wait for Clk_period;
		Addr <=  "00000000001111";
		Trees_din <= x"ff4f0095";
		wait for Clk_period;
		Addr <=  "00000000010000";
		Trees_din <= x"040b5208";
		wait for Clk_period;
		Addr <=  "00000000010001";
		Trees_din <= x"05045f04";
		wait for Clk_period;
		Addr <=  "00000000010010";
		Trees_din <= x"ff570095";
		wait for Clk_period;
		Addr <=  "00000000010011";
		Trees_din <= x"00270095";
		wait for Clk_period;
		Addr <=  "00000000010100";
		Trees_din <= x"01540095";
		wait for Clk_period;
		Addr <=  "00000000010101";
		Trees_din <= x"020d620c";
		wait for Clk_period;
		Addr <=  "00000000010110";
		Trees_din <= x"17004708";
		wait for Clk_period;
		Addr <=  "00000000010111";
		Trees_din <= x"01fc3604";
		wait for Clk_period;
		Addr <=  "00000000011000";
		Trees_din <= x"00b20095";
		wait for Clk_period;
		Addr <=  "00000000011001";
		Trees_din <= x"03590095";
		wait for Clk_period;
		Addr <=  "00000000011010";
		Trees_din <= x"00000095";
		wait for Clk_period;
		Addr <=  "00000000011011";
		Trees_din <= x"ff680095";
		wait for Clk_period;
		Addr <=  "00000000011100";
		Trees_din <= x"00c30f0c";
		wait for Clk_period;
		Addr <=  "00000000011101";
		Trees_din <= x"04171604";
		wait for Clk_period;
		Addr <=  "00000000011110";
		Trees_din <= x"ff530095";
		wait for Clk_period;
		Addr <=  "00000000011111";
		Trees_din <= x"00c00004";
		wait for Clk_period;
		Addr <=  "00000000100000";
		Trees_din <= x"ff6a0095";
		wait for Clk_period;
		Addr <=  "00000000100001";
		Trees_din <= x"02800095";
		wait for Clk_period;
		Addr <=  "00000000100010";
		Trees_din <= x"00d0a604";
		wait for Clk_period;
		Addr <=  "00000000100011";
		Trees_din <= x"01640095";
		wait for Clk_period;
		Addr <=  "00000000100100";
		Trees_din <= x"03b90095";
		wait for Clk_period;
		Addr <=  "00000000100101";
		Trees_din <= x"040ebb44";
		wait for Clk_period;
		Addr <=  "00000000100110";
		Trees_din <= x"0406af1c";
		wait for Clk_period;
		Addr <=  "00000000100111";
		Trees_din <= x"04048f0c";
		wait for Clk_period;
		Addr <=  "00000000101000";
		Trees_din <= x"1d013704";
		wait for Clk_period;
		Addr <=  "00000000101001";
		Trees_din <= x"ff550141";
		wait for Clk_period;
		Addr <=  "00000000101010";
		Trees_din <= x"0401f504";
		wait for Clk_period;
		Addr <=  "00000000101011";
		Trees_din <= x"ff730141";
		wait for Clk_period;
		Addr <=  "00000000101100";
		Trees_din <= x"00420141";
		wait for Clk_period;
		Addr <=  "00000000101101";
		Trees_din <= x"00f7bd04";
		wait for Clk_period;
		Addr <=  "00000000101110";
		Trees_din <= x"ff580141";
		wait for Clk_period;
		Addr <=  "00000000101111";
		Trees_din <= x"05fe0a08";
		wait for Clk_period;
		Addr <=  "00000000110000";
		Trees_din <= x"15053604";
		wait for Clk_period;
		Addr <=  "00000000110001";
		Trees_din <= x"ff790141";
		wait for Clk_period;
		Addr <=  "00000000110010";
		Trees_din <= x"002c0141";
		wait for Clk_period;
		Addr <=  "00000000110011";
		Trees_din <= x"011f0141";
		wait for Clk_period;
		Addr <=  "00000000110100";
		Trees_din <= x"00f01318";
		wait for Clk_period;
		Addr <=  "00000000110101";
		Trees_din <= x"00dc8808";
		wait for Clk_period;
		Addr <=  "00000000110110";
		Trees_din <= x"15f73a04";
		wait for Clk_period;
		Addr <=  "00000000110111";
		Trees_din <= x"001a0141";
		wait for Clk_period;
		Addr <=  "00000000111000";
		Trees_din <= x"ff560141";
		wait for Clk_period;
		Addr <=  "00000000111001";
		Trees_din <= x"05045f08";
		wait for Clk_period;
		Addr <=  "00000000111010";
		Trees_din <= x"13f7ac04";
		wait for Clk_period;
		Addr <=  "00000000111011";
		Trees_din <= x"00210141";
		wait for Clk_period;
		Addr <=  "00000000111100";
		Trees_din <= x"ff5f0141";
		wait for Clk_period;
		Addr <=  "00000000111101";
		Trees_din <= x"04081e04";
		wait for Clk_period;
		Addr <=  "00000000111110";
		Trees_din <= x"002c0141";
		wait for Clk_period;
		Addr <=  "00000000111111";
		Trees_din <= x"01670141";
		wait for Clk_period;
		Addr <=  "00000001000000";
		Trees_din <= x"02091208";
		wait for Clk_period;
		Addr <=  "00000001000001";
		Trees_din <= x"17004704";
		wait for Clk_period;
		Addr <=  "00000001000010";
		Trees_din <= x"01c00141";
		wait for Clk_period;
		Addr <=  "00000001000011";
		Trees_din <= x"000a0141";
		wait for Clk_period;
		Addr <=  "00000001000100";
		Trees_din <= x"0c020104";
		wait for Clk_period;
		Addr <=  "00000001000101";
		Trees_din <= x"ff730141";
		wait for Clk_period;
		Addr <=  "00000001000110";
		Trees_din <= x"00240141";
		wait for Clk_period;
		Addr <=  "00000001000111";
		Trees_din <= x"00c30f0c";
		wait for Clk_period;
		Addr <=  "00000001001000";
		Trees_din <= x"04171604";
		wait for Clk_period;
		Addr <=  "00000001001001";
		Trees_din <= x"ff5b0141";
		wait for Clk_period;
		Addr <=  "00000001001010";
		Trees_din <= x"00c00004";
		wait for Clk_period;
		Addr <=  "00000001001011";
		Trees_din <= x"ff730141";
		wait for Clk_period;
		Addr <=  "00000001001100";
		Trees_din <= x"01aa0141";
		wait for Clk_period;
		Addr <=  "00000001001101";
		Trees_din <= x"1103b804";
		wait for Clk_period;
		Addr <=  "00000001001110";
		Trees_din <= x"01af0141";
		wait for Clk_period;
		Addr <=  "00000001001111";
		Trees_din <= x"00880141";
		wait for Clk_period;
		Addr <=  "00000001010000";
		Trees_din <= x"040cd634";
		wait for Clk_period;
		Addr <=  "00000001010001";
		Trees_din <= x"04048f0c";
		wait for Clk_period;
		Addr <=  "00000001010010";
		Trees_din <= x"07003c08";
		wait for Clk_period;
		Addr <=  "00000001010011";
		Trees_din <= x"0fff1104";
		wait for Clk_period;
		Addr <=  "00000001010100";
		Trees_din <= x"003e01dd";
		wait for Clk_period;
		Addr <=  "00000001010101";
		Trees_din <= x"ff7b01dd";
		wait for Clk_period;
		Addr <=  "00000001010110";
		Trees_din <= x"ff5901dd";
		wait for Clk_period;
		Addr <=  "00000001010111";
		Trees_din <= x"00f01314";
		wait for Clk_period;
		Addr <=  "00000001011000";
		Trees_din <= x"0f04790c";
		wait for Clk_period;
		Addr <=  "00000001011001";
		Trees_din <= x"040bec04";
		wait for Clk_period;
		Addr <=  "00000001011010";
		Trees_din <= x"ff5a01dd";
		wait for Clk_period;
		Addr <=  "00000001011011";
		Trees_din <= x"0b026d04";
		wait for Clk_period;
		Addr <=  "00000001011100";
		Trees_din <= x"ff7b01dd";
		wait for Clk_period;
		Addr <=  "00000001011101";
		Trees_din <= x"003501dd";
		wait for Clk_period;
		Addr <=  "00000001011110";
		Trees_din <= x"1d00b804";
		wait for Clk_period;
		Addr <=  "00000001011111";
		Trees_din <= x"003601dd";
		wait for Clk_period;
		Addr <=  "00000001100000";
		Trees_din <= x"ff8001dd";
		wait for Clk_period;
		Addr <=  "00000001100001";
		Trees_din <= x"020d6210";
		wait for Clk_period;
		Addr <=  "00000001100010";
		Trees_din <= x"000a8008";
		wait for Clk_period;
		Addr <=  "00000001100011";
		Trees_din <= x"05f8b204";
		wait for Clk_period;
		Addr <=  "00000001100100";
		Trees_din <= x"ffa301dd";
		wait for Clk_period;
		Addr <=  "00000001100101";
		Trees_din <= x"013c01dd";
		wait for Clk_period;
		Addr <=  "00000001100110";
		Trees_din <= x"04078904";
		wait for Clk_period;
		Addr <=  "00000001100111";
		Trees_din <= x"ff6d01dd";
		wait for Clk_period;
		Addr <=  "00000001101000";
		Trees_din <= x"002701dd";
		wait for Clk_period;
		Addr <=  "00000001101001";
		Trees_din <= x"ff6701dd";
		wait for Clk_period;
		Addr <=  "00000001101010";
		Trees_din <= x"00c30f0c";
		wait for Clk_period;
		Addr <=  "00000001101011";
		Trees_din <= x"04171604";
		wait for Clk_period;
		Addr <=  "00000001101100";
		Trees_din <= x"ff5e01dd";
		wait for Clk_period;
		Addr <=  "00000001101101";
		Trees_din <= x"00c00004";
		wait for Clk_period;
		Addr <=  "00000001101110";
		Trees_din <= x"ff7a01dd";
		wait for Clk_period;
		Addr <=  "00000001101111";
		Trees_din <= x"014e01dd";
		wait for Clk_period;
		Addr <=  "00000001110000";
		Trees_din <= x"0116f10c";
		wait for Clk_period;
		Addr <=  "00000001110001";
		Trees_din <= x"0d038c04";
		wait for Clk_period;
		Addr <=  "00000001110010";
		Trees_din <= x"014901dd";
		wait for Clk_period;
		Addr <=  "00000001110011";
		Trees_din <= x"040fcf04";
		wait for Clk_period;
		Addr <=  "00000001110100";
		Trees_din <= x"ffa301dd";
		wait for Clk_period;
		Addr <=  "00000001110101";
		Trees_din <= x"00da01dd";
		wait for Clk_period;
		Addr <=  "00000001110110";
		Trees_din <= x"ff8701dd";
		wait for Clk_period;
		Addr <=  "00000001110111";
		Trees_din <= x"040cd634";
		wait for Clk_period;
		Addr <=  "00000001111000";
		Trees_din <= x"04048f0c";
		wait for Clk_period;
		Addr <=  "00000001111001";
		Trees_din <= x"1d013704";
		wait for Clk_period;
		Addr <=  "00000001111010";
		Trees_din <= x"ff5d0281";
		wait for Clk_period;
		Addr <=  "00000001111011";
		Trees_din <= x"14039904";
		wait for Clk_period;
		Addr <=  "00000001111100";
		Trees_din <= x"ff850281";
		wait for Clk_period;
		Addr <=  "00000001111101";
		Trees_din <= x"003a0281";
		wait for Clk_period;
		Addr <=  "00000001111110";
		Trees_din <= x"00f01314";
		wait for Clk_period;
		Addr <=  "00000001111111";
		Trees_din <= x"1603dc0c";
		wait for Clk_period;
		Addr <=  "00000010000000";
		Trees_din <= x"040bec04";
		wait for Clk_period;
		Addr <=  "00000010000001";
		Trees_din <= x"ff5e0281";
		wait for Clk_period;
		Addr <=  "00000010000010";
		Trees_din <= x"01096504";
		wait for Clk_period;
		Addr <=  "00000010000011";
		Trees_din <= x"00320281";
		wait for Clk_period;
		Addr <=  "00000010000100";
		Trees_din <= x"ff850281";
		wait for Clk_period;
		Addr <=  "00000010000101";
		Trees_din <= x"0d003704";
		wait for Clk_period;
		Addr <=  "00000010000110";
		Trees_din <= x"ff8b0281";
		wait for Clk_period;
		Addr <=  "00000010000111";
		Trees_din <= x"00360281";
		wait for Clk_period;
		Addr <=  "00000010001000";
		Trees_din <= x"020d6210";
		wait for Clk_period;
		Addr <=  "00000010001001";
		Trees_din <= x"000a8008";
		wait for Clk_period;
		Addr <=  "00000010001010";
		Trees_din <= x"05f8b204";
		wait for Clk_period;
		Addr <=  "00000010001011";
		Trees_din <= x"ffab0281";
		wait for Clk_period;
		Addr <=  "00000010001100";
		Trees_din <= x"00ea0281";
		wait for Clk_period;
		Addr <=  "00000010001101";
		Trees_din <= x"11004d04";
		wait for Clk_period;
		Addr <=  "00000010001110";
		Trees_din <= x"00310281";
		wait for Clk_period;
		Addr <=  "00000010001111";
		Trees_din <= x"ff720281";
		wait for Clk_period;
		Addr <=  "00000010010000";
		Trees_din <= x"ff6e0281";
		wait for Clk_period;
		Addr <=  "00000010010001";
		Trees_din <= x"00c30f0c";
		wait for Clk_period;
		Addr <=  "00000010010010";
		Trees_din <= x"04171604";
		wait for Clk_period;
		Addr <=  "00000010010011";
		Trees_din <= x"ff630281";
		wait for Clk_period;
		Addr <=  "00000010010100";
		Trees_din <= x"00c00004";
		wait for Clk_period;
		Addr <=  "00000010010101";
		Trees_din <= x"ff810281";
		wait for Clk_period;
		Addr <=  "00000010010110";
		Trees_din <= x"01180281";
		wait for Clk_period;
		Addr <=  "00000010010111";
		Trees_din <= x"0116f110";
		wait for Clk_period;
		Addr <=  "00000010011000";
		Trees_din <= x"020f190c";
		wait for Clk_period;
		Addr <=  "00000010011001";
		Trees_din <= x"0d03e008";
		wait for Clk_period;
		Addr <=  "00000010011010";
		Trees_din <= x"02fabf04";
		wait for Clk_period;
		Addr <=  "00000010011011";
		Trees_din <= x"00790281";
		wait for Clk_period;
		Addr <=  "00000010011100";
		Trees_din <= x"01190281";
		wait for Clk_period;
		Addr <=  "00000010011101";
		Trees_din <= x"00410281";
		wait for Clk_period;
		Addr <=  "00000010011110";
		Trees_din <= x"ffa40281";
		wait for Clk_period;
		Addr <=  "00000010011111";
		Trees_din <= x"ff920281";
		wait for Clk_period;
		Addr <=  "00000010100000";
		Trees_din <= x"040cd628";
		wait for Clk_period;
		Addr <=  "00000010100001";
		Trees_din <= x"04048f0c";
		wait for Clk_period;
		Addr <=  "00000010100010";
		Trees_din <= x"07003c08";
		wait for Clk_period;
		Addr <=  "00000010100011";
		Trees_din <= x"0904a304";
		wait for Clk_period;
		Addr <=  "00000010100100";
		Trees_din <= x"ff8e0315";
		wait for Clk_period;
		Addr <=  "00000010100101";
		Trees_din <= x"003b0315";
		wait for Clk_period;
		Addr <=  "00000010100110";
		Trees_din <= x"ff5f0315";
		wait for Clk_period;
		Addr <=  "00000010100111";
		Trees_din <= x"00f0130c";
		wait for Clk_period;
		Addr <=  "00000010101000";
		Trees_din <= x"0b038104";
		wait for Clk_period;
		Addr <=  "00000010101001";
		Trees_din <= x"ff610315";
		wait for Clk_period;
		Addr <=  "00000010101010";
		Trees_din <= x"16024b04";
		wait for Clk_period;
		Addr <=  "00000010101011";
		Trees_din <= x"ff730315";
		wait for Clk_period;
		Addr <=  "00000010101100";
		Trees_din <= x"00470315";
		wait for Clk_period;
		Addr <=  "00000010101101";
		Trees_din <= x"020d620c";
		wait for Clk_period;
		Addr <=  "00000010101110";
		Trees_din <= x"000fb808";
		wait for Clk_period;
		Addr <=  "00000010101111";
		Trees_din <= x"05f8e404";
		wait for Clk_period;
		Addr <=  "00000010110000";
		Trees_din <= x"ffa30315";
		wait for Clk_period;
		Addr <=  "00000010110001";
		Trees_din <= x"00b60315";
		wait for Clk_period;
		Addr <=  "00000010110010";
		Trees_din <= x"ff7c0315";
		wait for Clk_period;
		Addr <=  "00000010110011";
		Trees_din <= x"ff740315";
		wait for Clk_period;
		Addr <=  "00000010110100";
		Trees_din <= x"00c30f0c";
		wait for Clk_period;
		Addr <=  "00000010110101";
		Trees_din <= x"04171604";
		wait for Clk_period;
		Addr <=  "00000010110110";
		Trees_din <= x"ff670315";
		wait for Clk_period;
		Addr <=  "00000010110111";
		Trees_din <= x"00c00004";
		wait for Clk_period;
		Addr <=  "00000010111000";
		Trees_din <= x"ff880315";
		wait for Clk_period;
		Addr <=  "00000010111001";
		Trees_din <= x"00f60315";
		wait for Clk_period;
		Addr <=  "00000010111010";
		Trees_din <= x"0116f114";
		wait for Clk_period;
		Addr <=  "00000010111011";
		Trees_din <= x"07004d04";
		wait for Clk_period;
		Addr <=  "00000010111100";
		Trees_din <= x"00210315";
		wait for Clk_period;
		Addr <=  "00000010111101";
		Trees_din <= x"0d038c08";
		wait for Clk_period;
		Addr <=  "00000010111110";
		Trees_din <= x"09faf604";
		wait for Clk_period;
		Addr <=  "00000010111111";
		Trees_din <= x"008a0315";
		wait for Clk_period;
		Addr <=  "00000011000000";
		Trees_din <= x"00f50315";
		wait for Clk_period;
		Addr <=  "00000011000001";
		Trees_din <= x"19008b04";
		wait for Clk_period;
		Addr <=  "00000011000010";
		Trees_din <= x"00910315";
		wait for Clk_period;
		Addr <=  "00000011000011";
		Trees_din <= x"fffe0315";
		wait for Clk_period;
		Addr <=  "00000011000100";
		Trees_din <= x"ff9d0315";
		wait for Clk_period;
		Addr <=  "00000011000101";
		Trees_din <= x"040ac92c";
		wait for Clk_period;
		Addr <=  "00000011000110";
		Trees_din <= x"04048f0c";
		wait for Clk_period;
		Addr <=  "00000011000111";
		Trees_din <= x"1d013704";
		wait for Clk_period;
		Addr <=  "00000011001000";
		Trees_din <= x"ff6203a1";
		wait for Clk_period;
		Addr <=  "00000011001001";
		Trees_din <= x"1504e804";
		wait for Clk_period;
		Addr <=  "00000011001010";
		Trees_din <= x"ff9903a1";
		wait for Clk_period;
		Addr <=  "00000011001011";
		Trees_din <= x"003c03a1";
		wait for Clk_period;
		Addr <=  "00000011001100";
		Trees_din <= x"00f0130c";
		wait for Clk_period;
		Addr <=  "00000011001101";
		Trees_din <= x"0f047904";
		wait for Clk_period;
		Addr <=  "00000011001110";
		Trees_din <= x"ff6403a1";
		wait for Clk_period;
		Addr <=  "00000011001111";
		Trees_din <= x"11013104";
		wait for Clk_period;
		Addr <=  "00000011010000";
		Trees_din <= x"003803a1";
		wait for Clk_period;
		Addr <=  "00000011010001";
		Trees_din <= x"ffab03a1";
		wait for Clk_period;
		Addr <=  "00000011010010";
		Trees_din <= x"020d6210";
		wait for Clk_period;
		Addr <=  "00000011010011";
		Trees_din <= x"02ff3808";
		wait for Clk_period;
		Addr <=  "00000011010100";
		Trees_din <= x"02fa4c04";
		wait for Clk_period;
		Addr <=  "00000011010101";
		Trees_din <= x"003803a1";
		wait for Clk_period;
		Addr <=  "00000011010110";
		Trees_din <= x"ff6603a1";
		wait for Clk_period;
		Addr <=  "00000011010111";
		Trees_din <= x"000fb804";
		wait for Clk_period;
		Addr <=  "00000011011000";
		Trees_din <= x"009b03a1";
		wait for Clk_period;
		Addr <=  "00000011011001";
		Trees_din <= x"ffa603a1";
		wait for Clk_period;
		Addr <=  "00000011011010";
		Trees_din <= x"ff7c03a1";
		wait for Clk_period;
		Addr <=  "00000011011011";
		Trees_din <= x"00d0a614";
		wait for Clk_period;
		Addr <=  "00000011011100";
		Trees_din <= x"0417160c";
		wait for Clk_period;
		Addr <=  "00000011011101";
		Trees_din <= x"0c03b608";
		wait for Clk_period;
		Addr <=  "00000011011110";
		Trees_din <= x"09f72e04";
		wait for Clk_period;
		Addr <=  "00000011011111";
		Trees_din <= x"000703a1";
		wait for Clk_period;
		Addr <=  "00000011100000";
		Trees_din <= x"ff6603a1";
		wait for Clk_period;
		Addr <=  "00000011100001";
		Trees_din <= x"001203a1";
		wait for Clk_period;
		Addr <=  "00000011100010";
		Trees_din <= x"00c00004";
		wait for Clk_period;
		Addr <=  "00000011100011";
		Trees_din <= x"ff8f03a1";
		wait for Clk_period;
		Addr <=  "00000011100100";
		Trees_din <= x"00d903a1";
		wait for Clk_period;
		Addr <=  "00000011100101";
		Trees_din <= x"060e1c04";
		wait for Clk_period;
		Addr <=  "00000011100110";
		Trees_din <= x"00c303a1";
		wait for Clk_period;
		Addr <=  "00000011100111";
		Trees_din <= x"ffab03a1";
		wait for Clk_period;
		Addr <=  "00000011101000";
		Trees_din <= x"040ac934";
		wait for Clk_period;
		Addr <=  "00000011101001";
		Trees_din <= x"04048f0c";
		wait for Clk_period;
		Addr <=  "00000011101010";
		Trees_din <= x"07003c08";
		wait for Clk_period;
		Addr <=  "00000011101011";
		Trees_din <= x"0c015704";
		wait for Clk_period;
		Addr <=  "00000011101100";
		Trees_din <= x"00390445";
		wait for Clk_period;
		Addr <=  "00000011101101";
		Trees_din <= x"ffa30445";
		wait for Clk_period;
		Addr <=  "00000011101110";
		Trees_din <= x"ff640445";
		wait for Clk_period;
		Addr <=  "00000011101111";
		Trees_din <= x"00f1de0c";
		wait for Clk_period;
		Addr <=  "00000011110000";
		Trees_din <= x"1603dc08";
		wait for Clk_period;
		Addr <=  "00000011110001";
		Trees_din <= x"00f01304";
		wait for Clk_period;
		Addr <=  "00000011110010";
		Trees_din <= x"ff670445";
		wait for Clk_period;
		Addr <=  "00000011110011";
		Trees_din <= x"ffdc0445";
		wait for Clk_period;
		Addr <=  "00000011110100";
		Trees_din <= x"fff10445";
		wait for Clk_period;
		Addr <=  "00000011110101";
		Trees_din <= x"10021410";
		wait for Clk_period;
		Addr <=  "00000011110110";
		Trees_din <= x"04078908";
		wait for Clk_period;
		Addr <=  "00000011110111";
		Trees_din <= x"0ffd6404";
		wait for Clk_period;
		Addr <=  "00000011111000";
		Trees_din <= x"00030445";
		wait for Clk_period;
		Addr <=  "00000011111001";
		Trees_din <= x"ff650445";
		wait for Clk_period;
		Addr <=  "00000011111010";
		Trees_din <= x"19009f04";
		wait for Clk_period;
		Addr <=  "00000011111011";
		Trees_din <= x"ffdb0445";
		wait for Clk_period;
		Addr <=  "00000011111100";
		Trees_din <= x"00810445";
		wait for Clk_period;
		Addr <=  "00000011111101";
		Trees_din <= x"02088f08";
		wait for Clk_period;
		Addr <=  "00000011111110";
		Trees_din <= x"000fb804";
		wait for Clk_period;
		Addr <=  "00000011111111";
		Trees_din <= x"00e50445";
		wait for Clk_period;
		Addr <=  "00000100000000";
		Trees_din <= x"ffa70445";
		wait for Clk_period;
		Addr <=  "00000100000001";
		Trees_din <= x"ff950445";
		wait for Clk_period;
		Addr <=  "00000100000010";
		Trees_din <= x"00d0a60c";
		wait for Clk_period;
		Addr <=  "00000100000011";
		Trees_din <= x"04121004";
		wait for Clk_period;
		Addr <=  "00000100000100";
		Trees_din <= x"ff6b0445";
		wait for Clk_period;
		Addr <=  "00000100000101";
		Trees_din <= x"00c00004";
		wait for Clk_period;
		Addr <=  "00000100000110";
		Trees_din <= x"ff7c0445";
		wait for Clk_period;
		Addr <=  "00000100000111";
		Trees_din <= x"00b30445";
		wait for Clk_period;
		Addr <=  "00000100001000";
		Trees_din <= x"00d90008";
		wait for Clk_period;
		Addr <=  "00000100001001";
		Trees_din <= x"0c004e04";
		wait for Clk_period;
		Addr <=  "00000100001010";
		Trees_din <= x"009e0445";
		wait for Clk_period;
		Addr <=  "00000100001011";
		Trees_din <= x"ffc10445";
		wait for Clk_period;
		Addr <=  "00000100001100";
		Trees_din <= x"020b1e04";
		wait for Clk_period;
		Addr <=  "00000100001101";
		Trees_din <= x"00b90445";
		wait for Clk_period;
		Addr <=  "00000100001110";
		Trees_din <= x"1c003504";
		wait for Clk_period;
		Addr <=  "00000100001111";
		Trees_din <= x"ffed0445";
		wait for Clk_period;
		Addr <=  "00000100010000";
		Trees_din <= x"00860445";
		wait for Clk_period;
		Addr <=  "00000100010001";
		Trees_din <= x"040ac934";
		wait for Clk_period;
		Addr <=  "00000100010010";
		Trees_din <= x"04048f0c";
		wait for Clk_period;
		Addr <=  "00000100010011";
		Trees_din <= x"1d013704";
		wait for Clk_period;
		Addr <=  "00000100010100";
		Trees_din <= x"ff6504e1";
		wait for Clk_period;
		Addr <=  "00000100010101";
		Trees_din <= x"18002504";
		wait for Clk_period;
		Addr <=  "00000100010110";
		Trees_din <= x"ffb004e1";
		wait for Clk_period;
		Addr <=  "00000100010111";
		Trees_din <= x"003404e1";
		wait for Clk_period;
		Addr <=  "00000100011000";
		Trees_din <= x"00f1de0c";
		wait for Clk_period;
		Addr <=  "00000100011001";
		Trees_din <= x"0f047908";
		wait for Clk_period;
		Addr <=  "00000100011010";
		Trees_din <= x"00f01304";
		wait for Clk_period;
		Addr <=  "00000100011011";
		Trees_din <= x"ff6a04e1";
		wait for Clk_period;
		Addr <=  "00000100011100";
		Trees_din <= x"ffde04e1";
		wait for Clk_period;
		Addr <=  "00000100011101";
		Trees_din <= x"000004e1";
		wait for Clk_period;
		Addr <=  "00000100011110";
		Trees_din <= x"01fe8a0c";
		wait for Clk_period;
		Addr <=  "00000100011111";
		Trees_din <= x"03ff2308";
		wait for Clk_period;
		Addr <=  "00000100100000";
		Trees_din <= x"02091204";
		wait for Clk_period;
		Addr <=  "00000100100001";
		Trees_din <= x"004d04e1";
		wait for Clk_period;
		Addr <=  "00000100100010";
		Trees_din <= x"ffa904e1";
		wait for Clk_period;
		Addr <=  "00000100100011";
		Trees_din <= x"ff6c04e1";
		wait for Clk_period;
		Addr <=  "00000100100100";
		Trees_din <= x"03fc9208";
		wait for Clk_period;
		Addr <=  "00000100100101";
		Trees_din <= x"0efdce04";
		wait for Clk_period;
		Addr <=  "00000100100110";
		Trees_din <= x"fff304e1";
		wait for Clk_period;
		Addr <=  "00000100100111";
		Trees_din <= x"ff9b04e1";
		wait for Clk_period;
		Addr <=  "00000100101000";
		Trees_din <= x"09028804";
		wait for Clk_period;
		Addr <=  "00000100101001";
		Trees_din <= x"00ce04e1";
		wait for Clk_period;
		Addr <=  "00000100101010";
		Trees_din <= x"001e04e1";
		wait for Clk_period;
		Addr <=  "00000100101011";
		Trees_din <= x"00c30f0c";
		wait for Clk_period;
		Addr <=  "00000100101100";
		Trees_din <= x"04171604";
		wait for Clk_period;
		Addr <=  "00000100101101";
		Trees_din <= x"ff6f04e1";
		wait for Clk_period;
		Addr <=  "00000100101110";
		Trees_din <= x"00c00004";
		wait for Clk_period;
		Addr <=  "00000100101111";
		Trees_din <= x"ff9f04e1";
		wait for Clk_period;
		Addr <=  "00000100110000";
		Trees_din <= x"00ac04e1";
		wait for Clk_period;
		Addr <=  "00000100110001";
		Trees_din <= x"020f190c";
		wait for Clk_period;
		Addr <=  "00000100110010";
		Trees_din <= x"060e1c08";
		wait for Clk_period;
		Addr <=  "00000100110011";
		Trees_din <= x"0116f104";
		wait for Clk_period;
		Addr <=  "00000100110100";
		Trees_din <= x"00b904e1";
		wait for Clk_period;
		Addr <=  "00000100110101";
		Trees_din <= x"ffaa04e1";
		wait for Clk_period;
		Addr <=  "00000100110110";
		Trees_din <= x"ffa604e1";
		wait for Clk_period;
		Addr <=  "00000100110111";
		Trees_din <= x"ffa104e1";
		wait for Clk_period;
		Addr <=  "00000100111000";
		Trees_din <= x"0406af18";
		wait for Clk_period;
		Addr <=  "00000100111001";
		Trees_din <= x"02f6a804";
		wait for Clk_period;
		Addr <=  "00000100111010";
		Trees_din <= x"001c0545";
		wait for Clk_period;
		Addr <=  "00000100111011";
		Trees_din <= x"07003c04";
		wait for Clk_period;
		Addr <=  "00000100111100";
		Trees_din <= x"fff50545";
		wait for Clk_period;
		Addr <=  "00000100111101";
		Trees_din <= x"04034404";
		wait for Clk_period;
		Addr <=  "00000100111110";
		Trees_din <= x"ff660545";
		wait for Clk_period;
		Addr <=  "00000100111111";
		Trees_din <= x"04036104";
		wait for Clk_period;
		Addr <=  "00000101000000";
		Trees_din <= x"003c0545";
		wait for Clk_period;
		Addr <=  "00000101000001";
		Trees_din <= x"03fda304";
		wait for Clk_period;
		Addr <=  "00000101000010";
		Trees_din <= x"ffb70545";
		wait for Clk_period;
		Addr <=  "00000101000011";
		Trees_din <= x"ff6f0545";
		wait for Clk_period;
		Addr <=  "00000101000100";
		Trees_din <= x"020d6214";
		wait for Clk_period;
		Addr <=  "00000101000101";
		Trees_din <= x"06138010";
		wait for Clk_period;
		Addr <=  "00000101000110";
		Trees_din <= x"0118430c";
		wait for Clk_period;
		Addr <=  "00000101000111";
		Trees_din <= x"05109308";
		wait for Clk_period;
		Addr <=  "00000101001000";
		Trees_din <= x"040ac904";
		wait for Clk_period;
		Addr <=  "00000101001001";
		Trees_din <= x"004d0545";
		wait for Clk_period;
		Addr <=  "00000101001010";
		Trees_din <= x"00b10545";
		wait for Clk_period;
		Addr <=  "00000101001011";
		Trees_din <= x"ffb10545";
		wait for Clk_period;
		Addr <=  "00000101001100";
		Trees_din <= x"ff8d0545";
		wait for Clk_period;
		Addr <=  "00000101001101";
		Trees_din <= x"ff780545";
		wait for Clk_period;
		Addr <=  "00000101001110";
		Trees_din <= x"00f63204";
		wait for Clk_period;
		Addr <=  "00000101001111";
		Trees_din <= x"ff6e0545";
		wait for Clk_period;
		Addr <=  "00000101010000";
		Trees_din <= x"00000545";
		wait for Clk_period;
		Addr <=  "00000101010001";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00000101010010";
		Trees_din <= x"0406af18";
		wait for Clk_period;
		Addr <=  "00000101010011";
		Trees_din <= x"02f6a804";
		wait for Clk_period;
		Addr <=  "00000101010100";
		Trees_din <= x"002005b5";
		wait for Clk_period;
		Addr <=  "00000101010101";
		Trees_din <= x"1d013710";
		wait for Clk_period;
		Addr <=  "00000101010110";
		Trees_din <= x"04034404";
		wait for Clk_period;
		Addr <=  "00000101010111";
		Trees_din <= x"ff6705b5";
		wait for Clk_period;
		Addr <=  "00000101011000";
		Trees_din <= x"04036104";
		wait for Clk_period;
		Addr <=  "00000101011001";
		Trees_din <= x"003705b5";
		wait for Clk_period;
		Addr <=  "00000101011010";
		Trees_din <= x"15054204";
		wait for Clk_period;
		Addr <=  "00000101011011";
		Trees_din <= x"ff7e05b5";
		wait for Clk_period;
		Addr <=  "00000101011100";
		Trees_din <= x"ffe405b5";
		wait for Clk_period;
		Addr <=  "00000101011101";
		Trees_din <= x"000005b5";
		wait for Clk_period;
		Addr <=  "00000101011110";
		Trees_din <= x"020f191c";
		wait for Clk_period;
		Addr <=  "00000101011111";
		Trees_din <= x"060e1c14";
		wait for Clk_period;
		Addr <=  "00000101100000";
		Trees_din <= x"01184310";
		wait for Clk_period;
		Addr <=  "00000101100001";
		Trees_din <= x"0409a008";
		wait for Clk_period;
		Addr <=  "00000101100010";
		Trees_din <= x"00e76404";
		wait for Clk_period;
		Addr <=  "00000101100011";
		Trees_din <= x"ffa705b5";
		wait for Clk_period;
		Addr <=  "00000101100100";
		Trees_din <= x"006805b5";
		wait for Clk_period;
		Addr <=  "00000101100101";
		Trees_din <= x"0d039004";
		wait for Clk_period;
		Addr <=  "00000101100110";
		Trees_din <= x"00a505b5";
		wait for Clk_period;
		Addr <=  "00000101100111";
		Trees_din <= x"002505b5";
		wait for Clk_period;
		Addr <=  "00000101101000";
		Trees_din <= x"ff9405b5";
		wait for Clk_period;
		Addr <=  "00000101101001";
		Trees_din <= x"0c001a04";
		wait for Clk_period;
		Addr <=  "00000101101010";
		Trees_din <= x"001905b5";
		wait for Clk_period;
		Addr <=  "00000101101011";
		Trees_din <= x"ff7a05b5";
		wait for Clk_period;
		Addr <=  "00000101101100";
		Trees_din <= x"ff7305b5";
		wait for Clk_period;
		Addr <=  "00000101101101";
		Trees_din <= x"0406af18";
		wait for Clk_period;
		Addr <=  "00000101101110";
		Trees_din <= x"02f6a804";
		wait for Clk_period;
		Addr <=  "00000101101111";
		Trees_din <= x"00220619";
		wait for Clk_period;
		Addr <=  "00000101110000";
		Trees_din <= x"07003c04";
		wait for Clk_period;
		Addr <=  "00000101110001";
		Trees_din <= x"00050619";
		wait for Clk_period;
		Addr <=  "00000101110010";
		Trees_din <= x"04034404";
		wait for Clk_period;
		Addr <=  "00000101110011";
		Trees_din <= x"ff680619";
		wait for Clk_period;
		Addr <=  "00000101110100";
		Trees_din <= x"04036104";
		wait for Clk_period;
		Addr <=  "00000101110101";
		Trees_din <= x"00420619";
		wait for Clk_period;
		Addr <=  "00000101110110";
		Trees_din <= x"03fda304";
		wait for Clk_period;
		Addr <=  "00000101110111";
		Trees_din <= x"ffce0619";
		wait for Clk_period;
		Addr <=  "00000101111000";
		Trees_din <= x"ff770619";
		wait for Clk_period;
		Addr <=  "00000101111001";
		Trees_din <= x"020f1918";
		wait for Clk_period;
		Addr <=  "00000101111010";
		Trees_din <= x"06138014";
		wait for Clk_period;
		Addr <=  "00000101111011";
		Trees_din <= x"01184310";
		wait for Clk_period;
		Addr <=  "00000101111100";
		Trees_din <= x"040ac908";
		wait for Clk_period;
		Addr <=  "00000101111101";
		Trees_din <= x"00e76404";
		wait for Clk_period;
		Addr <=  "00000101111110";
		Trees_din <= x"ffa20619";
		wait for Clk_period;
		Addr <=  "00000101111111";
		Trees_din <= x"005b0619";
		wait for Clk_period;
		Addr <=  "00000110000000";
		Trees_din <= x"0d038c04";
		wait for Clk_period;
		Addr <=  "00000110000001";
		Trees_din <= x"009f0619";
		wait for Clk_period;
		Addr <=  "00000110000010";
		Trees_din <= x"00210619";
		wait for Clk_period;
		Addr <=  "00000110000011";
		Trees_din <= x"ff960619";
		wait for Clk_period;
		Addr <=  "00000110000100";
		Trees_din <= x"ff820619";
		wait for Clk_period;
		Addr <=  "00000110000101";
		Trees_din <= x"ff770619";
		wait for Clk_period;
		Addr <=  "00000110000110";
		Trees_din <= x"04048f18";
		wait for Clk_period;
		Addr <=  "00000110000111";
		Trees_din <= x"1d013714";
		wait for Clk_period;
		Addr <=  "00000110001000";
		Trees_din <= x"0403440c";
		wait for Clk_period;
		Addr <=  "00000110001001";
		Trees_din <= x"0b041c04";
		wait for Clk_period;
		Addr <=  "00000110001010";
		Trees_din <= x"ff67067d";
		wait for Clk_period;
		Addr <=  "00000110001011";
		Trees_din <= x"15fa8d04";
		wait for Clk_period;
		Addr <=  "00000110001100";
		Trees_din <= x"0048067d";
		wait for Clk_period;
		Addr <=  "00000110001101";
		Trees_din <= x"ff7f067d";
		wait for Clk_period;
		Addr <=  "00000110001110";
		Trees_din <= x"15f96504";
		wait for Clk_period;
		Addr <=  "00000110001111";
		Trees_din <= x"0041067d";
		wait for Clk_period;
		Addr <=  "00000110010000";
		Trees_din <= x"ff7f067d";
		wait for Clk_period;
		Addr <=  "00000110010001";
		Trees_din <= x"000d067d";
		wait for Clk_period;
		Addr <=  "00000110010010";
		Trees_din <= x"020f1918";
		wait for Clk_period;
		Addr <=  "00000110010011";
		Trees_din <= x"06138014";
		wait for Clk_period;
		Addr <=  "00000110010100";
		Trees_din <= x"0116f10c";
		wait for Clk_period;
		Addr <=  "00000110010101";
		Trees_din <= x"040b5208";
		wait for Clk_period;
		Addr <=  "00000110010110";
		Trees_din <= x"03017804";
		wait for Clk_period;
		Addr <=  "00000110010111";
		Trees_din <= x"003e067d";
		wait for Clk_period;
		Addr <=  "00000110011000";
		Trees_din <= x"ff78067d";
		wait for Clk_period;
		Addr <=  "00000110011001";
		Trees_din <= x"0095067d";
		wait for Clk_period;
		Addr <=  "00000110011010";
		Trees_din <= x"1200a004";
		wait for Clk_period;
		Addr <=  "00000110011011";
		Trees_din <= x"ff9c067d";
		wait for Clk_period;
		Addr <=  "00000110011100";
		Trees_din <= x"ffee067d";
		wait for Clk_period;
		Addr <=  "00000110011101";
		Trees_din <= x"ff84067d";
		wait for Clk_period;
		Addr <=  "00000110011110";
		Trees_din <= x"ff77067d";
		wait for Clk_period;
		Addr <=  "00000110011111";
		Trees_din <= x"04048f18";
		wait for Clk_period;
		Addr <=  "00000110100000";
		Trees_din <= x"07003c04";
		wait for Clk_period;
		Addr <=  "00000110100001";
		Trees_din <= x"001006e9";
		wait for Clk_period;
		Addr <=  "00000110100010";
		Trees_din <= x"0b041c0c";
		wait for Clk_period;
		Addr <=  "00000110100011";
		Trees_din <= x"04034404";
		wait for Clk_period;
		Addr <=  "00000110100100";
		Trees_din <= x"ff6806e9";
		wait for Clk_period;
		Addr <=  "00000110100101";
		Trees_din <= x"15f96504";
		wait for Clk_period;
		Addr <=  "00000110100110";
		Trees_din <= x"004506e9";
		wait for Clk_period;
		Addr <=  "00000110100111";
		Trees_din <= x"ff8806e9";
		wait for Clk_period;
		Addr <=  "00000110101000";
		Trees_din <= x"15fa8d04";
		wait for Clk_period;
		Addr <=  "00000110101001";
		Trees_din <= x"004806e9";
		wait for Clk_period;
		Addr <=  "00000110101010";
		Trees_din <= x"ff8406e9";
		wait for Clk_period;
		Addr <=  "00000110101011";
		Trees_din <= x"020f191c";
		wait for Clk_period;
		Addr <=  "00000110101100";
		Trees_din <= x"06138018";
		wait for Clk_period;
		Addr <=  "00000110101101";
		Trees_din <= x"040cd610";
		wait for Clk_period;
		Addr <=  "00000110101110";
		Trees_din <= x"03ffaf08";
		wait for Clk_period;
		Addr <=  "00000110101111";
		Trees_din <= x"010d0404";
		wait for Clk_period;
		Addr <=  "00000110110000";
		Trees_din <= x"005f06e9";
		wait for Clk_period;
		Addr <=  "00000110110001";
		Trees_din <= x"ffa406e9";
		wait for Clk_period;
		Addr <=  "00000110110010";
		Trees_din <= x"0a01a204";
		wait for Clk_period;
		Addr <=  "00000110110011";
		Trees_din <= x"ff7e06e9";
		wait for Clk_period;
		Addr <=  "00000110110100";
		Trees_din <= x"ffe906e9";
		wait for Clk_period;
		Addr <=  "00000110110101";
		Trees_din <= x"1c002c04";
		wait for Clk_period;
		Addr <=  "00000110110110";
		Trees_din <= x"002506e9";
		wait for Clk_period;
		Addr <=  "00000110110111";
		Trees_din <= x"007d06e9";
		wait for Clk_period;
		Addr <=  "00000110111000";
		Trees_din <= x"ff8a06e9";
		wait for Clk_period;
		Addr <=  "00000110111001";
		Trees_din <= x"ff7c06e9";
		wait for Clk_period;
		Addr <=  "00000110111010";
		Trees_din <= x"04048f18";
		wait for Clk_period;
		Addr <=  "00000110111011";
		Trees_din <= x"07003c04";
		wait for Clk_period;
		Addr <=  "00000110111100";
		Trees_din <= x"00100755";
		wait for Clk_period;
		Addr <=  "00000110111101";
		Trees_din <= x"0b041c0c";
		wait for Clk_period;
		Addr <=  "00000110111110";
		Trees_din <= x"04034404";
		wait for Clk_period;
		Addr <=  "00000110111111";
		Trees_din <= x"ff680755";
		wait for Clk_period;
		Addr <=  "00000111000000";
		Trees_din <= x"15f96b04";
		wait for Clk_period;
		Addr <=  "00000111000001";
		Trees_din <= x"00420755";
		wait for Clk_period;
		Addr <=  "00000111000010";
		Trees_din <= x"ff8f0755";
		wait for Clk_period;
		Addr <=  "00000111000011";
		Trees_din <= x"08005104";
		wait for Clk_period;
		Addr <=  "00000111000100";
		Trees_din <= x"004a0755";
		wait for Clk_period;
		Addr <=  "00000111000101";
		Trees_din <= x"ff8b0755";
		wait for Clk_period;
		Addr <=  "00000111000110";
		Trees_din <= x"020f191c";
		wait for Clk_period;
		Addr <=  "00000111000111";
		Trees_din <= x"06138018";
		wait for Clk_period;
		Addr <=  "00000111001000";
		Trees_din <= x"040ac90c";
		wait for Clk_period;
		Addr <=  "00000111001001";
		Trees_din <= x"03ffaf08";
		wait for Clk_period;
		Addr <=  "00000111001010";
		Trees_din <= x"010d0404";
		wait for Clk_period;
		Addr <=  "00000111001011";
		Trees_din <= x"004d0755";
		wait for Clk_period;
		Addr <=  "00000111001100";
		Trees_din <= x"ffac0755";
		wait for Clk_period;
		Addr <=  "00000111001101";
		Trees_din <= x"ff8d0755";
		wait for Clk_period;
		Addr <=  "00000111001110";
		Trees_din <= x"1100c804";
		wait for Clk_period;
		Addr <=  "00000111001111";
		Trees_din <= x"00120755";
		wait for Clk_period;
		Addr <=  "00000111010000";
		Trees_din <= x"020c5e04";
		wait for Clk_period;
		Addr <=  "00000111010001";
		Trees_din <= x"00770755";
		wait for Clk_period;
		Addr <=  "00000111010010";
		Trees_din <= x"001c0755";
		wait for Clk_period;
		Addr <=  "00000111010011";
		Trees_din <= x"ff920755";
		wait for Clk_period;
		Addr <=  "00000111010100";
		Trees_din <= x"ff810755";
		wait for Clk_period;
		Addr <=  "00000111010101";
		Trees_din <= x"04034410";
		wait for Clk_period;
		Addr <=  "00000111010110";
		Trees_din <= x"1c001e04";
		wait for Clk_period;
		Addr <=  "00000111010111";
		Trees_din <= x"000807b9";
		wait for Clk_period;
		Addr <=  "00000111011000";
		Trees_din <= x"0f046104";
		wait for Clk_period;
		Addr <=  "00000111011001";
		Trees_din <= x"ff6a07b9";
		wait for Clk_period;
		Addr <=  "00000111011010";
		Trees_din <= x"1d00d504";
		wait for Clk_period;
		Addr <=  "00000111011011";
		Trees_din <= x"ff9607b9";
		wait for Clk_period;
		Addr <=  "00000111011100";
		Trees_din <= x"004907b9";
		wait for Clk_period;
		Addr <=  "00000111011101";
		Trees_din <= x"020f1920";
		wait for Clk_period;
		Addr <=  "00000111011110";
		Trees_din <= x"03ffaf10";
		wait for Clk_period;
		Addr <=  "00000111011111";
		Trees_din <= x"0110ce0c";
		wait for Clk_period;
		Addr <=  "00000111100000";
		Trees_din <= x"000a8008";
		wait for Clk_period;
		Addr <=  "00000111100001";
		Trees_din <= x"0209d104";
		wait for Clk_period;
		Addr <=  "00000111100010";
		Trees_din <= x"008607b9";
		wait for Clk_period;
		Addr <=  "00000111100011";
		Trees_din <= x"000707b9";
		wait for Clk_period;
		Addr <=  "00000111100100";
		Trees_din <= x"ffd907b9";
		wait for Clk_period;
		Addr <=  "00000111100101";
		Trees_din <= x"ffc907b9";
		wait for Clk_period;
		Addr <=  "00000111100110";
		Trees_din <= x"040ac904";
		wait for Clk_period;
		Addr <=  "00000111100111";
		Trees_din <= x"ff8107b9";
		wait for Clk_period;
		Addr <=  "00000111101000";
		Trees_din <= x"04121008";
		wait for Clk_period;
		Addr <=  "00000111101001";
		Trees_din <= x"00d0a604";
		wait for Clk_period;
		Addr <=  "00000111101010";
		Trees_din <= x"ffa707b9";
		wait for Clk_period;
		Addr <=  "00000111101011";
		Trees_din <= x"004407b9";
		wait for Clk_period;
		Addr <=  "00000111101100";
		Trees_din <= x"005707b9";
		wait for Clk_period;
		Addr <=  "00000111101101";
		Trees_din <= x"ff8407b9";
		wait for Clk_period;
		Addr <=  "00000111101110";
		Trees_din <= x"04034410";
		wait for Clk_period;
		Addr <=  "00000111101111";
		Trees_din <= x"0b041c08";
		wait for Clk_period;
		Addr <=  "00000111110000";
		Trees_din <= x"1a003004";
		wait for Clk_period;
		Addr <=  "00000111110001";
		Trees_din <= x"fffb0835";
		wait for Clk_period;
		Addr <=  "00000111110010";
		Trees_din <= x"ff6b0835";
		wait for Clk_period;
		Addr <=  "00000111110011";
		Trees_din <= x"02fcdf04";
		wait for Clk_period;
		Addr <=  "00000111110100";
		Trees_din <= x"00480835";
		wait for Clk_period;
		Addr <=  "00000111110101";
		Trees_din <= x"ffa10835";
		wait for Clk_period;
		Addr <=  "00000111110110";
		Trees_din <= x"020f192c";
		wait for Clk_period;
		Addr <=  "00000111110111";
		Trees_din <= x"03ffaf1c";
		wait for Clk_period;
		Addr <=  "00000111111000";
		Trees_din <= x"1d00c410";
		wait for Clk_period;
		Addr <=  "00000111111001";
		Trees_din <= x"05fc6c08";
		wait for Clk_period;
		Addr <=  "00000111111010";
		Trees_din <= x"03fdf304";
		wait for Clk_period;
		Addr <=  "00000111111011";
		Trees_din <= x"ffb20835";
		wait for Clk_period;
		Addr <=  "00000111111100";
		Trees_din <= x"ffec0835";
		wait for Clk_period;
		Addr <=  "00000111111101";
		Trees_din <= x"1b019e04";
		wait for Clk_period;
		Addr <=  "00000111111110";
		Trees_din <= x"00030835";
		wait for Clk_period;
		Addr <=  "00000111111111";
		Trees_din <= x"00420835";
		wait for Clk_period;
		Addr <=  "00001000000000";
		Trees_din <= x"17003c04";
		wait for Clk_period;
		Addr <=  "00001000000001";
		Trees_din <= x"fffb0835";
		wait for Clk_period;
		Addr <=  "00001000000010";
		Trees_din <= x"19009904";
		wait for Clk_period;
		Addr <=  "00001000000011";
		Trees_din <= x"00200835";
		wait for Clk_period;
		Addr <=  "00001000000100";
		Trees_din <= x"009f0835";
		wait for Clk_period;
		Addr <=  "00001000000101";
		Trees_din <= x"040cd608";
		wait for Clk_period;
		Addr <=  "00001000000110";
		Trees_din <= x"03017804";
		wait for Clk_period;
		Addr <=  "00001000000111";
		Trees_din <= x"ffcf0835";
		wait for Clk_period;
		Addr <=  "00001000001000";
		Trees_din <= x"ff820835";
		wait for Clk_period;
		Addr <=  "00001000001001";
		Trees_din <= x"04121004";
		wait for Clk_period;
		Addr <=  "00001000001010";
		Trees_din <= x"00010835";
		wait for Clk_period;
		Addr <=  "00001000001011";
		Trees_din <= x"004f0835";
		wait for Clk_period;
		Addr <=  "00001000001100";
		Trees_din <= x"ff8a0835";
		wait for Clk_period;
		Addr <=  "00001000001101";
		Trees_din <= x"04034410";
		wait for Clk_period;
		Addr <=  "00001000001110";
		Trees_din <= x"0f046108";
		wait for Clk_period;
		Addr <=  "00001000001111";
		Trees_din <= x"1a003004";
		wait for Clk_period;
		Addr <=  "00001000010000";
		Trees_din <= x"fffc0891";
		wait for Clk_period;
		Addr <=  "00001000010001";
		Trees_din <= x"ff6c0891";
		wait for Clk_period;
		Addr <=  "00001000010010";
		Trees_din <= x"1b024504";
		wait for Clk_period;
		Addr <=  "00001000010011";
		Trees_din <= x"ffac0891";
		wait for Clk_period;
		Addr <=  "00001000010100";
		Trees_din <= x"004a0891";
		wait for Clk_period;
		Addr <=  "00001000010101";
		Trees_din <= x"020f191c";
		wait for Clk_period;
		Addr <=  "00001000010110";
		Trees_din <= x"02ff0f08";
		wait for Clk_period;
		Addr <=  "00001000010111";
		Trees_din <= x"01ffcd04";
		wait for Clk_period;
		Addr <=  "00001000011000";
		Trees_din <= x"ff8d0891";
		wait for Clk_period;
		Addr <=  "00001000011001";
		Trees_din <= x"00170891";
		wait for Clk_period;
		Addr <=  "00001000011010";
		Trees_din <= x"0109650c";
		wait for Clk_period;
		Addr <=  "00001000011011";
		Trees_din <= x"02097e08";
		wait for Clk_period;
		Addr <=  "00001000011100";
		Trees_din <= x"1d00da04";
		wait for Clk_period;
		Addr <=  "00001000011101";
		Trees_din <= x"00760891";
		wait for Clk_period;
		Addr <=  "00001000011110";
		Trees_din <= x"00020891";
		wait for Clk_period;
		Addr <=  "00001000011111";
		Trees_din <= x"fff90891";
		wait for Clk_period;
		Addr <=  "00001000100000";
		Trees_din <= x"04121004";
		wait for Clk_period;
		Addr <=  "00001000100001";
		Trees_din <= x"ffa40891";
		wait for Clk_period;
		Addr <=  "00001000100010";
		Trees_din <= x"00520891";
		wait for Clk_period;
		Addr <=  "00001000100011";
		Trees_din <= x"ff910891";
		wait for Clk_period;
		Addr <=  "00001000100100";
		Trees_din <= x"0406af1c";
		wait for Clk_period;
		Addr <=  "00001000100101";
		Trees_din <= x"0b041c14";
		wait for Clk_period;
		Addr <=  "00001000100110";
		Trees_din <= x"04029c04";
		wait for Clk_period;
		Addr <=  "00001000100111";
		Trees_din <= x"ff6e08f5";
		wait for Clk_period;
		Addr <=  "00001000101000";
		Trees_din <= x"16028808";
		wait for Clk_period;
		Addr <=  "00001000101001";
		Trees_din <= x"1900a204";
		wait for Clk_period;
		Addr <=  "00001000101010";
		Trees_din <= x"ff8008f5";
		wait for Clk_period;
		Addr <=  "00001000101011";
		Trees_din <= x"ffe108f5";
		wait for Clk_period;
		Addr <=  "00001000101100";
		Trees_din <= x"09050404";
		wait for Clk_period;
		Addr <=  "00001000101101";
		Trees_din <= x"ffd408f5";
		wait for Clk_period;
		Addr <=  "00001000101110";
		Trees_din <= x"006008f5";
		wait for Clk_period;
		Addr <=  "00001000101111";
		Trees_din <= x"02fb8e04";
		wait for Clk_period;
		Addr <=  "00001000110000";
		Trees_din <= x"009808f5";
		wait for Clk_period;
		Addr <=  "00001000110001";
		Trees_din <= x"ffa208f5";
		wait for Clk_period;
		Addr <=  "00001000110010";
		Trees_din <= x"00d9000c";
		wait for Clk_period;
		Addr <=  "00001000110011";
		Trees_din <= x"04171608";
		wait for Clk_period;
		Addr <=  "00001000110100";
		Trees_din <= x"00d0a604";
		wait for Clk_period;
		Addr <=  "00001000110101";
		Trees_din <= x"ffa208f5";
		wait for Clk_period;
		Addr <=  "00001000110110";
		Trees_din <= x"fff908f5";
		wait for Clk_period;
		Addr <=  "00001000110111";
		Trees_din <= x"003108f5";
		wait for Clk_period;
		Addr <=  "00001000111000";
		Trees_din <= x"01fe0a04";
		wait for Clk_period;
		Addr <=  "00001000111001";
		Trees_din <= x"fff308f5";
		wait for Clk_period;
		Addr <=  "00001000111010";
		Trees_din <= x"19009e04";
		wait for Clk_period;
		Addr <=  "00001000111011";
		Trees_din <= x"006608f5";
		wait for Clk_period;
		Addr <=  "00001000111100";
		Trees_din <= x"001608f5";
		wait for Clk_period;
		Addr <=  "00001000111101";
		Trees_din <= x"04014b04";
		wait for Clk_period;
		Addr <=  "00001000111110";
		Trees_din <= x"ff720949";
		wait for Clk_period;
		Addr <=  "00001000111111";
		Trees_din <= x"000fb824";
		wait for Clk_period;
		Addr <=  "00001001000000";
		Trees_din <= x"00fcab18";
		wait for Clk_period;
		Addr <=  "00001001000001";
		Trees_din <= x"040cd60c";
		wait for Clk_period;
		Addr <=  "00001001000010";
		Trees_din <= x"1100a708";
		wait for Clk_period;
		Addr <=  "00001001000011";
		Trees_din <= x"03fe5204";
		wait for Clk_period;
		Addr <=  "00001001000100";
		Trees_din <= x"00160949";
		wait for Clk_period;
		Addr <=  "00001001000101";
		Trees_din <= x"ffd60949";
		wait for Clk_period;
		Addr <=  "00001001000110";
		Trees_din <= x"ff940949";
		wait for Clk_period;
		Addr <=  "00001001000111";
		Trees_din <= x"020bd208";
		wait for Clk_period;
		Addr <=  "00001001001000";
		Trees_din <= x"05fe8204";
		wait for Clk_period;
		Addr <=  "00001001001001";
		Trees_din <= x"00110949";
		wait for Clk_period;
		Addr <=  "00001001001010";
		Trees_din <= x"00550949";
		wait for Clk_period;
		Addr <=  "00001001001011";
		Trees_din <= x"ffe50949";
		wait for Clk_period;
		Addr <=  "00001001001100";
		Trees_din <= x"1a004508";
		wait for Clk_period;
		Addr <=  "00001001001101";
		Trees_din <= x"18003804";
		wait for Clk_period;
		Addr <=  "00001001001110";
		Trees_din <= x"00420949";
		wait for Clk_period;
		Addr <=  "00001001001111";
		Trees_din <= x"00ec0949";
		wait for Clk_period;
		Addr <=  "00001001010000";
		Trees_din <= x"ffdf0949";
		wait for Clk_period;
		Addr <=  "00001001010001";
		Trees_din <= x"ff830949";
		wait for Clk_period;
		Addr <=  "00001001010010";
		Trees_din <= x"04014b04";
		wait for Clk_period;
		Addr <=  "00001001010011";
		Trees_din <= x"ff750995";
		wait for Clk_period;
		Addr <=  "00001001010100";
		Trees_din <= x"000fb820";
		wait for Clk_period;
		Addr <=  "00001001010101";
		Trees_din <= x"00fcab14";
		wait for Clk_period;
		Addr <=  "00001001010110";
		Trees_din <= x"040ac908";
		wait for Clk_period;
		Addr <=  "00001001010111";
		Trees_din <= x"1100a704";
		wait for Clk_period;
		Addr <=  "00001001011000";
		Trees_din <= x"fffd0995";
		wait for Clk_period;
		Addr <=  "00001001011001";
		Trees_din <= x"ff890995";
		wait for Clk_period;
		Addr <=  "00001001011010";
		Trees_din <= x"020bd208";
		wait for Clk_period;
		Addr <=  "00001001011011";
		Trees_din <= x"04121004";
		wait for Clk_period;
		Addr <=  "00001001011100";
		Trees_din <= x"00160995";
		wait for Clk_period;
		Addr <=  "00001001011101";
		Trees_din <= x"00560995";
		wait for Clk_period;
		Addr <=  "00001001011110";
		Trees_din <= x"ffe30995";
		wait for Clk_period;
		Addr <=  "00001001011111";
		Trees_din <= x"1a004508";
		wait for Clk_period;
		Addr <=  "00001001100000";
		Trees_din <= x"05fe0104";
		wait for Clk_period;
		Addr <=  "00001001100001";
		Trees_din <= x"00290995";
		wait for Clk_period;
		Addr <=  "00001001100010";
		Trees_din <= x"00c70995";
		wait for Clk_period;
		Addr <=  "00001001100011";
		Trees_din <= x"ffe20995";
		wait for Clk_period;
		Addr <=  "00001001100100";
		Trees_din <= x"ff8a0995";
		wait for Clk_period;
		Addr <=  "00001001100101";
		Trees_din <= x"04014b04";
		wait for Clk_period;
		Addr <=  "00001001100110";
		Trees_din <= x"ff7909e1";
		wait for Clk_period;
		Addr <=  "00001001100111";
		Trees_din <= x"000fb820";
		wait for Clk_period;
		Addr <=  "00001001101000";
		Trees_din <= x"0003dc18";
		wait for Clk_period;
		Addr <=  "00001001101001";
		Trees_din <= x"040ac90c";
		wait for Clk_period;
		Addr <=  "00001001101010";
		Trees_din <= x"10028708";
		wait for Clk_period;
		Addr <=  "00001001101011";
		Trees_din <= x"05fba004";
		wait for Clk_period;
		Addr <=  "00001001101100";
		Trees_din <= x"ffe209e1";
		wait for Clk_period;
		Addr <=  "00001001101101";
		Trees_din <= x"ff9009e1";
		wait for Clk_period;
		Addr <=  "00001001101110";
		Trees_din <= x"000c09e1";
		wait for Clk_period;
		Addr <=  "00001001101111";
		Trees_din <= x"00d0a608";
		wait for Clk_period;
		Addr <=  "00001001110000";
		Trees_din <= x"08005704";
		wait for Clk_period;
		Addr <=  "00001001110001";
		Trees_din <= x"ffc809e1";
		wait for Clk_period;
		Addr <=  "00001001110010";
		Trees_din <= x"001009e1";
		wait for Clk_period;
		Addr <=  "00001001110011";
		Trees_din <= x"005909e1";
		wait for Clk_period;
		Addr <=  "00001001110100";
		Trees_din <= x"10022204";
		wait for Clk_period;
		Addr <=  "00001001110101";
		Trees_din <= x"000109e1";
		wait for Clk_period;
		Addr <=  "00001001110110";
		Trees_din <= x"00a609e1";
		wait for Clk_period;
		Addr <=  "00001001110111";
		Trees_din <= x"ff9109e1";
		wait for Clk_period;
		Addr <=  "00001001111000";
		Trees_din <= x"04014b04";
		wait for Clk_period;
		Addr <=  "00001001111001";
		Trees_din <= x"ff7d0a1d";
		wait for Clk_period;
		Addr <=  "00001001111010";
		Trees_din <= x"0f046118";
		wait for Clk_period;
		Addr <=  "00001001111011";
		Trees_din <= x"04078908";
		wait for Clk_period;
		Addr <=  "00001001111100";
		Trees_din <= x"16028804";
		wait for Clk_period;
		Addr <=  "00001001111101";
		Trees_din <= x"ff950a1d";
		wait for Clk_period;
		Addr <=  "00001001111110";
		Trees_din <= x"00030a1d";
		wait for Clk_period;
		Addr <=  "00001001111111";
		Trees_din <= x"0116f10c";
		wait for Clk_period;
		Addr <=  "00001010000000";
		Trees_din <= x"16000004";
		wait for Clk_period;
		Addr <=  "00001010000001";
		Trees_din <= x"ffe20a1d";
		wait for Clk_period;
		Addr <=  "00001010000010";
		Trees_din <= x"03012c04";
		wait for Clk_period;
		Addr <=  "00001010000011";
		Trees_din <= x"00630a1d";
		wait for Clk_period;
		Addr <=  "00001010000100";
		Trees_din <= x"00140a1d";
		wait for Clk_period;
		Addr <=  "00001010000101";
		Trees_din <= x"ffc20a1d";
		wait for Clk_period;
		Addr <=  "00001010000110";
		Trees_din <= x"00690a1d";
		wait for Clk_period;
		Addr <=  "00001010000111";
		Trees_din <= x"04014b04";
		wait for Clk_period;
		Addr <=  "00001010001000";
		Trees_din <= x"ff820a59";
		wait for Clk_period;
		Addr <=  "00001010001001";
		Trees_din <= x"03ff0110";
		wait for Clk_period;
		Addr <=  "00001010001010";
		Trees_din <= x"1d00c508";
		wait for Clk_period;
		Addr <=  "00001010001011";
		Trees_din <= x"00f7bd04";
		wait for Clk_period;
		Addr <=  "00001010001100";
		Trees_din <= x"00040a59";
		wait for Clk_period;
		Addr <=  "00001010001101";
		Trees_din <= x"ffc00a59";
		wait for Clk_period;
		Addr <=  "00001010001110";
		Trees_din <= x"17003e04";
		wait for Clk_period;
		Addr <=  "00001010001111";
		Trees_din <= x"ffff0a59";
		wait for Clk_period;
		Addr <=  "00001010010000";
		Trees_din <= x"00840a59";
		wait for Clk_period;
		Addr <=  "00001010010001";
		Trees_din <= x"040ebb08";
		wait for Clk_period;
		Addr <=  "00001010010010";
		Trees_din <= x"11030104";
		wait for Clk_period;
		Addr <=  "00001010010011";
		Trees_din <= x"ff9a0a59";
		wait for Clk_period;
		Addr <=  "00001010010100";
		Trees_din <= x"ffeb0a59";
		wait for Clk_period;
		Addr <=  "00001010010101";
		Trees_din <= x"00210a59";
		wait for Clk_period;
		Addr <=  "00001010010110";
		Trees_din <= x"04014b04";
		wait for Clk_period;
		Addr <=  "00001010010111";
		Trees_din <= x"ff870a8d";
		wait for Clk_period;
		Addr <=  "00001010011000";
		Trees_din <= x"0f046114";
		wait for Clk_period;
		Addr <=  "00001010011001";
		Trees_din <= x"04078908";
		wait for Clk_period;
		Addr <=  "00001010011010";
		Trees_din <= x"16028804";
		wait for Clk_period;
		Addr <=  "00001010011011";
		Trees_din <= x"ff9f0a8d";
		wait for Clk_period;
		Addr <=  "00001010011100";
		Trees_din <= x"00020a8d";
		wait for Clk_period;
		Addr <=  "00001010011101";
		Trees_din <= x"00d90008";
		wait for Clk_period;
		Addr <=  "00001010011110";
		Trees_din <= x"1b022404";
		wait for Clk_period;
		Addr <=  "00001010011111";
		Trees_din <= x"ffd20a8d";
		wait for Clk_period;
		Addr <=  "00001010100000";
		Trees_din <= x"00070a8d";
		wait for Clk_period;
		Addr <=  "00001010100001";
		Trees_din <= x"00460a8d";
		wait for Clk_period;
		Addr <=  "00001010100010";
		Trees_din <= x"00590a8d";
		wait for Clk_period;
		Addr <=  "00001010100011";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00001010100100";
		Trees_din <= x"04014b04";
		wait for Clk_period;
		Addr <=  "00001010100101";
		Trees_din <= x"ff8c0ac5";
		wait for Clk_period;
		Addr <=  "00001010100110";
		Trees_din <= x"03ff120c";
		wait for Clk_period;
		Addr <=  "00001010100111";
		Trees_din <= x"1d00c504";
		wait for Clk_period;
		Addr <=  "00001010101000";
		Trees_din <= x"ffdc0ac5";
		wait for Clk_period;
		Addr <=  "00001010101001";
		Trees_din <= x"17003e04";
		wait for Clk_period;
		Addr <=  "00001010101010";
		Trees_din <= x"00020ac5";
		wait for Clk_period;
		Addr <=  "00001010101011";
		Trees_din <= x"00730ac5";
		wait for Clk_period;
		Addr <=  "00001010101100";
		Trees_din <= x"040ac904";
		wait for Clk_period;
		Addr <=  "00001010101101";
		Trees_din <= x"ffa90ac5";
		wait for Clk_period;
		Addr <=  "00001010101110";
		Trees_din <= x"1b02cf04";
		wait for Clk_period;
		Addr <=  "00001010101111";
		Trees_din <= x"fff40ac5";
		wait for Clk_period;
		Addr <=  "00001010110000";
		Trees_din <= x"00290ac5";
		wait for Clk_period;
		Addr <=  "00001010110001";
		Trees_din <= x"04014b04";
		wait for Clk_period;
		Addr <=  "00001010110010";
		Trees_din <= x"ff910af9";
		wait for Clk_period;
		Addr <=  "00001010110011";
		Trees_din <= x"03ff380c";
		wait for Clk_period;
		Addr <=  "00001010110100";
		Trees_din <= x"1d00c504";
		wait for Clk_period;
		Addr <=  "00001010110101";
		Trees_din <= x"ffe00af9";
		wait for Clk_period;
		Addr <=  "00001010110110";
		Trees_din <= x"12009804";
		wait for Clk_period;
		Addr <=  "00001010110111";
		Trees_din <= x"00700af9";
		wait for Clk_period;
		Addr <=  "00001010111000";
		Trees_din <= x"000c0af9";
		wait for Clk_period;
		Addr <=  "00001010111001";
		Trees_din <= x"040ebb08";
		wait for Clk_period;
		Addr <=  "00001010111010";
		Trees_din <= x"0c00cc04";
		wait for Clk_period;
		Addr <=  "00001010111011";
		Trees_din <= x"ffe60af9";
		wait for Clk_period;
		Addr <=  "00001010111100";
		Trees_din <= x"ffa60af9";
		wait for Clk_period;
		Addr <=  "00001010111101";
		Trees_din <= x"001b0af9";
		wait for Clk_period;
		Addr <=  "00001010111110";
		Trees_din <= x"04014b04";
		wait for Clk_period;
		Addr <=  "00001010111111";
		Trees_din <= x"ff960b2d";
		wait for Clk_period;
		Addr <=  "00001011000000";
		Trees_din <= x"0f046114";
		wait for Clk_period;
		Addr <=  "00001011000001";
		Trees_din <= x"04078908";
		wait for Clk_period;
		Addr <=  "00001011000010";
		Trees_din <= x"16028804";
		wait for Clk_period;
		Addr <=  "00001011000011";
		Trees_din <= x"ffac0b2d";
		wait for Clk_period;
		Addr <=  "00001011000100";
		Trees_din <= x"00010b2d";
		wait for Clk_period;
		Addr <=  "00001011000101";
		Trees_din <= x"00d90008";
		wait for Clk_period;
		Addr <=  "00001011000110";
		Trees_din <= x"12009204";
		wait for Clk_period;
		Addr <=  "00001011000111";
		Trees_din <= x"00030b2d";
		wait for Clk_period;
		Addr <=  "00001011001000";
		Trees_din <= x"ffe30b2d";
		wait for Clk_period;
		Addr <=  "00001011001001";
		Trees_din <= x"00410b2d";
		wait for Clk_period;
		Addr <=  "00001011001010";
		Trees_din <= x"00470b2d";
		wait for Clk_period;
		Addr <=  "00001011001011";
		Trees_din <= x"04014b04";
		wait for Clk_period;
		Addr <=  "00001011001100";
		Trees_din <= x"ff9c0b61";
		wait for Clk_period;
		Addr <=  "00001011001101";
		Trees_din <= x"03ff380c";
		wait for Clk_period;
		Addr <=  "00001011001110";
		Trees_din <= x"18003a08";
		wait for Clk_period;
		Addr <=  "00001011001111";
		Trees_din <= x"10020004";
		wait for Clk_period;
		Addr <=  "00001011010000";
		Trees_din <= x"fffd0b61";
		wait for Clk_period;
		Addr <=  "00001011010001";
		Trees_din <= x"005f0b61";
		wait for Clk_period;
		Addr <=  "00001011010010";
		Trees_din <= x"ffdf0b61";
		wait for Clk_period;
		Addr <=  "00001011010011";
		Trees_din <= x"040fcf08";
		wait for Clk_period;
		Addr <=  "00001011010100";
		Trees_din <= x"0c00cc04";
		wait for Clk_period;
		Addr <=  "00001011010101";
		Trees_din <= x"ffea0b61";
		wait for Clk_period;
		Addr <=  "00001011010110";
		Trees_din <= x"ffb10b61";
		wait for Clk_period;
		Addr <=  "00001011010111";
		Trees_din <= x"001b0b61";
		wait for Clk_period;
		Addr <=  "00001011011000";
		Trees_din <= x"04014b04";
		wait for Clk_period;
		Addr <=  "00001011011001";
		Trees_din <= x"ffa10b8d";
		wait for Clk_period;
		Addr <=  "00001011011010";
		Trees_din <= x"0f046110";
		wait for Clk_period;
		Addr <=  "00001011011011";
		Trees_din <= x"04078908";
		wait for Clk_period;
		Addr <=  "00001011011100";
		Trees_din <= x"10022d04";
		wait for Clk_period;
		Addr <=  "00001011011101";
		Trees_din <= x"ffb00b8d";
		wait for Clk_period;
		Addr <=  "00001011011110";
		Trees_din <= x"fffa0b8d";
		wait for Clk_period;
		Addr <=  "00001011011111";
		Trees_din <= x"020a6904";
		wait for Clk_period;
		Addr <=  "00001011100000";
		Trees_din <= x"00340b8d";
		wait for Clk_period;
		Addr <=  "00001011100001";
		Trees_din <= x"ffea0b8d";
		wait for Clk_period;
		Addr <=  "00001011100010";
		Trees_din <= x"003c0b8d";
		wait for Clk_period;
		Addr <=  "00001011100011";
		Trees_din <= x"04014b04";
		wait for Clk_period;
		Addr <=  "00001011100100";
		Trees_din <= x"ffa60bb9";
		wait for Clk_period;
		Addr <=  "00001011100101";
		Trees_din <= x"03ff380c";
		wait for Clk_period;
		Addr <=  "00001011100110";
		Trees_din <= x"1d00c504";
		wait for Clk_period;
		Addr <=  "00001011100111";
		Trees_din <= x"ffe40bb9";
		wait for Clk_period;
		Addr <=  "00001011101000";
		Trees_din <= x"12009804";
		wait for Clk_period;
		Addr <=  "00001011101001";
		Trees_din <= x"00590bb9";
		wait for Clk_period;
		Addr <=  "00001011101010";
		Trees_din <= x"00060bb9";
		wait for Clk_period;
		Addr <=  "00001011101011";
		Trees_din <= x"040ac904";
		wait for Clk_period;
		Addr <=  "00001011101100";
		Trees_din <= x"ffbc0bb9";
		wait for Clk_period;
		Addr <=  "00001011101101";
		Trees_din <= x"000e0bb9";
		wait for Clk_period;
		Addr <=  "00001011101110";
		Trees_din <= x"0406af08";
		wait for Clk_period;
		Addr <=  "00001011101111";
		Trees_din <= x"08005104";
		wait for Clk_period;
		Addr <=  "00001011110000";
		Trees_din <= x"00190bd5";
		wait for Clk_period;
		Addr <=  "00001011110001";
		Trees_din <= x"ffa30bd5";
		wait for Clk_period;
		Addr <=  "00001011110010";
		Trees_din <= x"00d90004";
		wait for Clk_period;
		Addr <=  "00001011110011";
		Trees_din <= x"ffeb0bd5";
		wait for Clk_period;
		Addr <=  "00001011110100";
		Trees_din <= x"00350bd5";
		wait for Clk_period;
		Addr <=  "00001011110101";
		Trees_din <= x"04014b04";
		wait for Clk_period;
		Addr <=  "00001011110110";
		Trees_din <= x"ffae0c01";
		wait for Clk_period;
		Addr <=  "00001011110111";
		Trees_din <= x"020a6910";
		wait for Clk_period;
		Addr <=  "00001011111000";
		Trees_din <= x"03ff1208";
		wait for Clk_period;
		Addr <=  "00001011111001";
		Trees_din <= x"10023f04";
		wait for Clk_period;
		Addr <=  "00001011111010";
		Trees_din <= x"fffb0c01";
		wait for Clk_period;
		Addr <=  "00001011111011";
		Trees_din <= x"004d0c01";
		wait for Clk_period;
		Addr <=  "00001011111100";
		Trees_din <= x"02019004";
		wait for Clk_period;
		Addr <=  "00001011111101";
		Trees_din <= x"ffd40c01";
		wait for Clk_period;
		Addr <=  "00001011111110";
		Trees_din <= x"00150c01";
		wait for Clk_period;
		Addr <=  "00001011111111";
		Trees_din <= x"ffda0c01";
		wait for Clk_period;
		Addr <=  "00001100000000";
		Trees_din <= x"0406af08";
		wait for Clk_period;
		Addr <=  "00001100000001";
		Trees_din <= x"08005104";
		wait for Clk_period;
		Addr <=  "00001100000010";
		Trees_din <= x"00140c1d";
		wait for Clk_period;
		Addr <=  "00001100000011";
		Trees_din <= x"ffaa0c1d";
		wait for Clk_period;
		Addr <=  "00001100000100";
		Trees_din <= x"00d90004";
		wait for Clk_period;
		Addr <=  "00001100000101";
		Trees_din <= x"fff10c1d";
		wait for Clk_period;
		Addr <=  "00001100000110";
		Trees_din <= x"00300c1d";
		wait for Clk_period;
		Addr <=  "00001100000111";
		Trees_din <= x"040db70c";
		wait for Clk_period;
		Addr <=  "00001100001000";
		Trees_din <= x"10022d04";
		wait for Clk_period;
		Addr <=  "00001100001001";
		Trees_din <= x"ffbf0c39";
		wait for Clk_period;
		Addr <=  "00001100001010";
		Trees_din <= x"13fc3704";
		wait for Clk_period;
		Addr <=  "00001100001011";
		Trees_din <= x"00330c39";
		wait for Clk_period;
		Addr <=  "00001100001100";
		Trees_din <= x"ffdf0c39";
		wait for Clk_period;
		Addr <=  "00001100001101";
		Trees_din <= x"00270c39";
		wait for Clk_period;
		Addr <=  "00001100001110";
		Trees_din <= x"0406af08";
		wait for Clk_period;
		Addr <=  "00001100001111";
		Trees_din <= x"08005104";
		wait for Clk_period;
		Addr <=  "00001100010000";
		Trees_din <= x"00100c55";
		wait for Clk_period;
		Addr <=  "00001100010001";
		Trees_din <= x"ffb30c55";
		wait for Clk_period;
		Addr <=  "00001100010010";
		Trees_din <= x"020a6904";
		wait for Clk_period;
		Addr <=  "00001100010011";
		Trees_din <= x"00280c55";
		wait for Clk_period;
		Addr <=  "00001100010100";
		Trees_din <= x"fff20c55";
		wait for Clk_period;
		Addr <=  "00001100010101";
		Trees_din <= x"04073408";
		wait for Clk_period;
		Addr <=  "00001100010110";
		Trees_din <= x"0effd004";
		wait for Clk_period;
		Addr <=  "00001100010111";
		Trees_din <= x"ffb70c71";
		wait for Clk_period;
		Addr <=  "00001100011000";
		Trees_din <= x"00080c71";
		wait for Clk_period;
		Addr <=  "00001100011001";
		Trees_din <= x"00d90004";
		wait for Clk_period;
		Addr <=  "00001100011010";
		Trees_din <= x"fff20c71";
		wait for Clk_period;
		Addr <=  "00001100011011";
		Trees_din <= x"002f0c71";
		wait for Clk_period;
		Addr <=  "00001100011100";
		Trees_din <= x"040db70c";
		wait for Clk_period;
		Addr <=  "00001100011101";
		Trees_din <= x"1a004508";
		wait for Clk_period;
		Addr <=  "00001100011110";
		Trees_din <= x"12009804";
		wait for Clk_period;
		Addr <=  "00001100011111";
		Trees_din <= x"00360c8d";
		wait for Clk_period;
		Addr <=  "00001100100000";
		Trees_din <= x"ffd40c8d";
		wait for Clk_period;
		Addr <=  "00001100100001";
		Trees_din <= x"ffc20c8d";
		wait for Clk_period;
		Addr <=  "00001100100010";
		Trees_din <= x"00240c8d";
		wait for Clk_period;
		Addr <=  "00001100100011";
		Trees_din <= x"0406af08";
		wait for Clk_period;
		Addr <=  "00001100100100";
		Trees_din <= x"08005104";
		wait for Clk_period;
		Addr <=  "00001100100101";
		Trees_din <= x"000e0ca9";
		wait for Clk_period;
		Addr <=  "00001100100110";
		Trees_din <= x"ffbd0ca9";
		wait for Clk_period;
		Addr <=  "00001100100111";
		Trees_din <= x"00d90004";
		wait for Clk_period;
		Addr <=  "00001100101000";
		Trees_din <= x"fff20ca9";
		wait for Clk_period;
		Addr <=  "00001100101001";
		Trees_din <= x"002b0ca9";
		wait for Clk_period;
		Addr <=  "00001100101010";
		Trees_din <= x"040cd60c";
		wait for Clk_period;
		Addr <=  "00001100101011";
		Trees_din <= x"10022d04";
		wait for Clk_period;
		Addr <=  "00001100101100";
		Trees_din <= x"ffc70cc5";
		wait for Clk_period;
		Addr <=  "00001100101101";
		Trees_din <= x"0a01e504";
		wait for Clk_period;
		Addr <=  "00001100101110";
		Trees_din <= x"fffd0cc5";
		wait for Clk_period;
		Addr <=  "00001100101111";
		Trees_din <= x"00120cc5";
		wait for Clk_period;
		Addr <=  "00001100110000";
		Trees_din <= x"00200cc5";
		wait for Clk_period;
		Addr <=  "00001100110001";
		Trees_din <= x"04073408";
		wait for Clk_period;
		Addr <=  "00001100110010";
		Trees_din <= x"0effd004";
		wait for Clk_period;
		Addr <=  "00001100110011";
		Trees_din <= x"ffc30ce1";
		wait for Clk_period;
		Addr <=  "00001100110100";
		Trees_din <= x"00080ce1";
		wait for Clk_period;
		Addr <=  "00001100110101";
		Trees_din <= x"0d01ca04";
		wait for Clk_period;
		Addr <=  "00001100110110";
		Trees_din <= x"00270ce1";
		wait for Clk_period;
		Addr <=  "00001100110111";
		Trees_din <= x"fff40ce1";
		wait for Clk_period;
		Addr <=  "00001100111000";
		Trees_din <= x"04073408";
		wait for Clk_period;
		Addr <=  "00001100111001";
		Trees_din <= x"17004004";
		wait for Clk_period;
		Addr <=  "00001100111010";
		Trees_din <= x"00070cfd";
		wait for Clk_period;
		Addr <=  "00001100111011";
		Trees_din <= x"ffc40cfd";
		wait for Clk_period;
		Addr <=  "00001100111100";
		Trees_din <= x"00dc8804";
		wait for Clk_period;
		Addr <=  "00001100111101";
		Trees_din <= x"fff40cfd";
		wait for Clk_period;
		Addr <=  "00001100111110";
		Trees_din <= x"002c0cfd";
		wait for Clk_period;
		Addr <=  "00001100111111";
		Trees_din <= x"040db708";
		wait for Clk_period;
		Addr <=  "00001101000000";
		Trees_din <= x"10022d04";
		wait for Clk_period;
		Addr <=  "00001101000001";
		Trees_din <= x"ffd00d11";
		wait for Clk_period;
		Addr <=  "00001101000010";
		Trees_din <= x"00090d11";
		wait for Clk_period;
		Addr <=  "00001101000011";
		Trees_din <= x"001f0d11";
		wait for Clk_period;
		Addr <=  "00001101000100";
		Trees_din <= x"0406af08";
		wait for Clk_period;
		Addr <=  "00001101000101";
		Trees_din <= x"07005504";
		wait for Clk_period;
		Addr <=  "00001101000110";
		Trees_din <= x"00070d2d";
		wait for Clk_period;
		Addr <=  "00001101000111";
		Trees_din <= x"ffc70d2d";
		wait for Clk_period;
		Addr <=  "00001101001000";
		Trees_din <= x"12009304";
		wait for Clk_period;
		Addr <=  "00001101001001";
		Trees_din <= x"00240d2d";
		wait for Clk_period;
		Addr <=  "00001101001010";
		Trees_din <= x"fff80d2d";
		wait for Clk_period;
		Addr <=  "00001101001011";
		Trees_din <= x"0406af08";
		wait for Clk_period;
		Addr <=  "00001101001100";
		Trees_din <= x"0effd304";
		wait for Clk_period;
		Addr <=  "00001101001101";
		Trees_din <= x"ffce0d49";
		wait for Clk_period;
		Addr <=  "00001101001110";
		Trees_din <= x"00040d49";
		wait for Clk_period;
		Addr <=  "00001101001111";
		Trees_din <= x"03ff8e04";
		wait for Clk_period;
		Addr <=  "00001101010000";
		Trees_din <= x"00230d49";
		wait for Clk_period;
		Addr <=  "00001101010001";
		Trees_din <= x"fff90d49";
		wait for Clk_period;
		Addr <=  "00001101010010";
		Trees_din <= x"040cd60c";
		wait for Clk_period;
		Addr <=  "00001101010011";
		Trees_din <= x"1a004508";
		wait for Clk_period;
		Addr <=  "00001101010100";
		Trees_din <= x"06fed504";
		wait for Clk_period;
		Addr <=  "00001101010101";
		Trees_din <= x"001e0d65";
		wait for Clk_period;
		Addr <=  "00001101010110";
		Trees_din <= x"ffee0d65";
		wait for Clk_period;
		Addr <=  "00001101010111";
		Trees_din <= x"ffcd0d65";
		wait for Clk_period;
		Addr <=  "00001101011000";
		Trees_din <= x"001a0d65";
		wait for Clk_period;
		Addr <=  "00001101011001";
		Trees_din <= x"04073408";
		wait for Clk_period;
		Addr <=  "00001101011010";
		Trees_din <= x"0effd004";
		wait for Clk_period;
		Addr <=  "00001101011011";
		Trees_din <= x"ffcf0d81";
		wait for Clk_period;
		Addr <=  "00001101011100";
		Trees_din <= x"00060d81";
		wait for Clk_period;
		Addr <=  "00001101011101";
		Trees_din <= x"12009304";
		wait for Clk_period;
		Addr <=  "00001101011110";
		Trees_din <= x"00220d81";
		wait for Clk_period;
		Addr <=  "00001101011111";
		Trees_din <= x"fff70d81";
		wait for Clk_period;
		Addr <=  "00001101100000";
		Trees_din <= x"16000104";
		wait for Clk_period;
		Addr <=  "00001101100001";
		Trees_din <= x"ffde0d9d";
		wait for Clk_period;
		Addr <=  "00001101100010";
		Trees_din <= x"01069b08";
		wait for Clk_period;
		Addr <=  "00001101100011";
		Trees_din <= x"13fc7c04";
		wait for Clk_period;
		Addr <=  "00001101100100";
		Trees_din <= x"00200d9d";
		wait for Clk_period;
		Addr <=  "00001101100101";
		Trees_din <= x"00070d9d";
		wait for Clk_period;
		Addr <=  "00001101100110";
		Trees_din <= x"ffee0d9d";
		wait for Clk_period;
		Addr <=  "00001101100111";
		Trees_din <= x"0406af04";
		wait for Clk_period;
		Addr <=  "00001101101000";
		Trees_din <= x"ffe40db1";
		wait for Clk_period;
		Addr <=  "00001101101001";
		Trees_din <= x"03ff8e04";
		wait for Clk_period;
		Addr <=  "00001101101010";
		Trees_din <= x"00220db1";
		wait for Clk_period;
		Addr <=  "00001101101011";
		Trees_din <= x"fffa0db1";
		wait for Clk_period;
		Addr <=  "00001101101100";
		Trees_din <= x"16000104";
		wait for Clk_period;
		Addr <=  "00001101101101";
		Trees_din <= x"ffe10dc5";
		wait for Clk_period;
		Addr <=  "00001101101110";
		Trees_din <= x"0405a904";
		wait for Clk_period;
		Addr <=  "00001101101111";
		Trees_din <= x"fff10dc5";
		wait for Clk_period;
		Addr <=  "00001101110000";
		Trees_din <= x"001b0dc5";
		wait for Clk_period;
		Addr <=  "00001101110001";
		Trees_din <= x"12009808";
		wait for Clk_period;
		Addr <=  "00001101110010";
		Trees_din <= x"18003a04";
		wait for Clk_period;
		Addr <=  "00001101110011";
		Trees_din <= x"002b0dd9";
		wait for Clk_period;
		Addr <=  "00001101110100";
		Trees_din <= x"ffeb0dd9";
		wait for Clk_period;
		Addr <=  "00001101110101";
		Trees_din <= x"ffe60dd9";
		wait for Clk_period;
		Addr <=  "00001101110110";
		Trees_din <= x"040cd608";
		wait for Clk_period;
		Addr <=  "00001101110111";
		Trees_din <= x"02ffbf04";
		wait for Clk_period;
		Addr <=  "00001101111000";
		Trees_din <= x"000e0ded";
		wait for Clk_period;
		Addr <=  "00001101111001";
		Trees_din <= x"ffd80ded";
		wait for Clk_period;
		Addr <=  "00001101111010";
		Trees_din <= x"00190ded";
		wait for Clk_period;
		Addr <=  "00001101111011";
		Trees_din <= x"04048f04";
		wait for Clk_period;
		Addr <=  "00001101111100";
		Trees_din <= x"ffe30e01";
		wait for Clk_period;
		Addr <=  "00001101111101";
		Trees_din <= x"00f01304";
		wait for Clk_period;
		Addr <=  "00001101111110";
		Trees_din <= x"fff50e01";
		wait for Clk_period;
		Addr <=  "00001101111111";
		Trees_din <= x"00240e01";
		wait for Clk_period;
		Addr <=  "00001110000000";
		Trees_din <= x"18003a08";
		wait for Clk_period;
		Addr <=  "00001110000001";
		Trees_din <= x"18003704";
		wait for Clk_period;
		Addr <=  "00001110000010";
		Trees_din <= x"ffef0e15";
		wait for Clk_period;
		Addr <=  "00001110000011";
		Trees_din <= x"00270e15";
		wait for Clk_period;
		Addr <=  "00001110000100";
		Trees_din <= x"ffea0e15";
		wait for Clk_period;
		Addr <=  "00001110000101";
		Trees_din <= x"040cd608";
		wait for Clk_period;
		Addr <=  "00001110000110";
		Trees_din <= x"10022d04";
		wait for Clk_period;
		Addr <=  "00001110000111";
		Trees_din <= x"ffd80e29";
		wait for Clk_period;
		Addr <=  "00001110001000";
		Trees_din <= x"00080e29";
		wait for Clk_period;
		Addr <=  "00001110001001";
		Trees_din <= x"001a0e29";
		wait for Clk_period;
		Addr <=  "00001110001010";
		Trees_din <= x"0406af04";
		wait for Clk_period;
		Addr <=  "00001110001011";
		Trees_din <= x"ffe80e3d";
		wait for Clk_period;
		Addr <=  "00001110001100";
		Trees_din <= x"12009304";
		wait for Clk_period;
		Addr <=  "00001110001101";
		Trees_din <= x"001e0e3d";
		wait for Clk_period;
		Addr <=  "00001110001110";
		Trees_din <= x"fffc0e3d";
		wait for Clk_period;
		Addr <=  "00001110001111";
		Trees_din <= x"18003a08";
		wait for Clk_period;
		Addr <=  "00001110010000";
		Trees_din <= x"12009804";
		wait for Clk_period;
		Addr <=  "00001110010001";
		Trees_din <= x"00250e51";
		wait for Clk_period;
		Addr <=  "00001110010010";
		Trees_din <= x"fff00e51";
		wait for Clk_period;
		Addr <=  "00001110010011";
		Trees_din <= x"ffea0e51";
		wait for Clk_period;
		Addr <=  "00001110010100";
		Trees_din <= x"03ffaf08";
		wait for Clk_period;
		Addr <=  "00001110010101";
		Trees_din <= x"03fdd404";
		wait for Clk_period;
		Addr <=  "00001110010110";
		Trees_din <= x"ffee0e65";
		wait for Clk_period;
		Addr <=  "00001110010111";
		Trees_din <= x"00240e65";
		wait for Clk_period;
		Addr <=  "00001110011000";
		Trees_din <= x"ffeb0e65";
		wait for Clk_period;
		Addr <=  "00001110011001";
		Trees_din <= x"05001708";
		wait for Clk_period;
		Addr <=  "00001110011010";
		Trees_din <= x"14027804";
		wait for Clk_period;
		Addr <=  "00001110011011";
		Trees_din <= x"00040e79";
		wait for Clk_period;
		Addr <=  "00001110011100";
		Trees_din <= x"000f0e79";
		wait for Clk_period;
		Addr <=  "00001110011101";
		Trees_din <= x"ffec0e79";
		wait for Clk_period;
		Addr <=  "00001110011110";
		Trees_din <= x"040cd608";
		wait for Clk_period;
		Addr <=  "00001110011111";
		Trees_din <= x"1d00d004";
		wait for Clk_period;
		Addr <=  "00001110100000";
		Trees_din <= x"ffdc0e8d";
		wait for Clk_period;
		Addr <=  "00001110100001";
		Trees_din <= x"00070e8d";
		wait for Clk_period;
		Addr <=  "00001110100010";
		Trees_din <= x"00190e8d";
		wait for Clk_period;
		Addr <=  "00001110100011";
		Trees_din <= x"04048f04";
		wait for Clk_period;
		Addr <=  "00001110100100";
		Trees_din <= x"ffe50ea1";
		wait for Clk_period;
		Addr <=  "00001110100101";
		Trees_din <= x"00f01304";
		wait for Clk_period;
		Addr <=  "00001110100110";
		Trees_din <= x"fff70ea1";
		wait for Clk_period;
		Addr <=  "00001110100111";
		Trees_din <= x"00220ea1";
		wait for Clk_period;
		Addr <=  "00001110101000";
		Trees_din <= x"040cd608";
		wait for Clk_period;
		Addr <=  "00001110101001";
		Trees_din <= x"00fcab04";
		wait for Clk_period;
		Addr <=  "00001110101010";
		Trees_din <= x"ffdc0eb5";
		wait for Clk_period;
		Addr <=  "00001110101011";
		Trees_din <= x"00070eb5";
		wait for Clk_period;
		Addr <=  "00001110101100";
		Trees_din <= x"00180eb5";
		wait for Clk_period;
		Addr <=  "00001110101101";
		Trees_din <= x"0406af04";
		wait for Clk_period;
		Addr <=  "00001110101110";
		Trees_din <= x"ffe90ec1";
		wait for Clk_period;
		Addr <=  "00001110101111";
		Trees_din <= x"00110ec1";
		wait for Clk_period;
		Addr <=  "00001110110000";
		Trees_din <= x"03ffaf08";
		wait for Clk_period;
		Addr <=  "00001110110001";
		Trees_din <= x"03fdd404";
		wait for Clk_period;
		Addr <=  "00001110110010";
		Trees_din <= x"fff10ed5";
		wait for Clk_period;
		Addr <=  "00001110110011";
		Trees_din <= x"00200ed5";
		wait for Clk_period;
		Addr <=  "00001110110100";
		Trees_din <= x"ffeb0ed5";
		wait for Clk_period;
		Addr <=  "00001110110101";
		Trees_din <= x"18003a04";
		wait for Clk_period;
		Addr <=  "00001110110110";
		Trees_din <= x"000b0ee1";
		wait for Clk_period;
		Addr <=  "00001110110111";
		Trees_din <= x"ffed0ee1";
		wait for Clk_period;
		Addr <=  "00001110111000";
		Trees_din <= x"19008f04";
		wait for Clk_period;
		Addr <=  "00001110111001";
		Trees_din <= x"000f0ef5";
		wait for Clk_period;
		Addr <=  "00001110111010";
		Trees_din <= x"0d015804";
		wait for Clk_period;
		Addr <=  "00001110111011";
		Trees_din <= x"00090ef5";
		wait for Clk_period;
		Addr <=  "00001110111100";
		Trees_din <= x"ffe10ef5";
		wait for Clk_period;
		Addr <=  "00001110111101";
		Trees_din <= x"05001704";
		wait for Clk_period;
		Addr <=  "00001110111110";
		Trees_din <= x"000c0f01";
		wait for Clk_period;
		Addr <=  "00001110111111";
		Trees_din <= x"ffee0f01";
		wait for Clk_period;
		Addr <=  "00001111000000";
		Trees_din <= x"18003a04";
		wait for Clk_period;
		Addr <=  "00001111000001";
		Trees_din <= x"000b0f0d";
		wait for Clk_period;
		Addr <=  "00001111000010";
		Trees_din <= x"ffee0f0d";
		wait for Clk_period;
		Addr <=  "00001111000011";
		Trees_din <= x"0efd6f04";
		wait for Clk_period;
		Addr <=  "00001111000100";
		Trees_din <= x"000f0f21";
		wait for Clk_period;
		Addr <=  "00001111000101";
		Trees_din <= x"0a015904";
		wait for Clk_period;
		Addr <=  "00001111000110";
		Trees_din <= x"ffe20f21";
		wait for Clk_period;
		Addr <=  "00001111000111";
		Trees_din <= x"000b0f21";
		wait for Clk_period;
		Addr <=  "00001111001000";
		Trees_din <= x"12009804";
		wait for Clk_period;
		Addr <=  "00001111001001";
		Trees_din <= x"000a0f2d";
		wait for Clk_period;
		Addr <=  "00001111001010";
		Trees_din <= x"ffee0f2d";
		wait for Clk_period;
		Addr <=  "00001111001011";
		Trees_din <= x"05ffe604";
		wait for Clk_period;
		Addr <=  "00001111001100";
		Trees_din <= x"000b0f39";
		wait for Clk_period;
		Addr <=  "00001111001101";
		Trees_din <= x"fff00f39";
		wait for Clk_period;
		Addr <=  "00001111001110";
		Trees_din <= x"0efd6f04";
		wait for Clk_period;
		Addr <=  "00001111001111";
		Trees_din <= x"000f0f4d";
		wait for Clk_period;
		Addr <=  "00001111010000";
		Trees_din <= x"1b022404";
		wait for Clk_period;
		Addr <=  "00001111010001";
		Trees_din <= x"ffea0f4d";
		wait for Clk_period;
		Addr <=  "00001111010010";
		Trees_din <= x"00020f4d";
		wait for Clk_period;
		Addr <=  "00001111010011";
		Trees_din <= x"03ffaf04";
		wait for Clk_period;
		Addr <=  "00001111010100";
		Trees_din <= x"000a0f59";
		wait for Clk_period;
		Addr <=  "00001111010101";
		Trees_din <= x"ffef0f59";
		wait for Clk_period;
		Addr <=  "00001111010110";
		Trees_din <= x"15028604";
		wait for Clk_period;
		Addr <=  "00001111010111";
		Trees_din <= x"fff10f65";
		wait for Clk_period;
		Addr <=  "00001111011000";
		Trees_din <= x"000b0f65";
		wait for Clk_period;
		Addr <=  "00001111011001";
		Trees_din <= x"05001704";
		wait for Clk_period;
		Addr <=  "00001111011010";
		Trees_din <= x"000a0f71";
		wait for Clk_period;
		Addr <=  "00001111011011";
		Trees_din <= x"fff00f71";
		wait for Clk_period;
		Addr <=  "00001111011100";
		Trees_din <= x"18003a04";
		wait for Clk_period;
		Addr <=  "00001111011101";
		Trees_din <= x"00090f7d";
		wait for Clk_period;
		Addr <=  "00001111011110";
		Trees_din <= x"fff00f7d";
		wait for Clk_period;
		Addr <=  "00001111011111";
		Trees_din <= x"19008f04";
		wait for Clk_period;
		Addr <=  "00001111100000";
		Trees_din <= x"000d0f89";
		wait for Clk_period;
		Addr <=  "00001111100001";
		Trees_din <= x"fff30f89";
		wait for Clk_period;
		Addr <=  "00001111100010";
		Trees_din <= x"18003a04";
		wait for Clk_period;
		Addr <=  "00001111100011";
		Trees_din <= x"00090f95";
		wait for Clk_period;
		Addr <=  "00001111100100";
		Trees_din <= x"fff10f95";
		wait for Clk_period;
		Addr <=  "00001111100101";
		Trees_din <= x"19008f04";
		wait for Clk_period;
		Addr <=  "00001111100110";
		Trees_din <= x"000d0fa1";
		wait for Clk_period;
		Addr <=  "00001111100111";
		Trees_din <= x"fff40fa1";
		wait for Clk_period;
		Addr <=  "00001111101000";
		Trees_din <= x"16006904";
		wait for Clk_period;
		Addr <=  "00001111101001";
		Trees_din <= x"fff30fad";
		wait for Clk_period;
		Addr <=  "00001111101010";
		Trees_din <= x"000b0fad";
		wait for Clk_period;
		Addr <=  "00001111101011";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  6
        -----------
		Addr <=  "00000000000000";
		Trees_din <= x"030faf14";
		wait for Clk_period;
		Addr <=  "00000000000001";
		Trees_din <= x"030b980c";
		wait for Clk_period;
		Addr <=  "00000000000010";
		Trees_din <= x"03092d04";
		wait for Clk_period;
		Addr <=  "00000000000011";
		Trees_din <= x"ff4d0035";
		wait for Clk_period;
		Addr <=  "00000000000100";
		Trees_din <= x"00f0ae04";
		wait for Clk_period;
		Addr <=  "00000000000101";
		Trees_din <= x"ff590035";
		wait for Clk_period;
		Addr <=  "00000000000110";
		Trees_din <= x"02500035";
		wait for Clk_period;
		Addr <=  "00000000000111";
		Trees_din <= x"00e9ab04";
		wait for Clk_period;
		Addr <=  "00000000001000";
		Trees_din <= x"ff5d0035";
		wait for Clk_period;
		Addr <=  "00000000001001";
		Trees_din <= x"03840035";
		wait for Clk_period;
		Addr <=  "00000000001010";
		Trees_din <= x"06138004";
		wait for Clk_period;
		Addr <=  "00000000001011";
		Trees_din <= x"03e50035";
		wait for Clk_period;
		Addr <=  "00000000001100";
		Trees_din <= x"ff7d0035";
		wait for Clk_period;
		Addr <=  "00000000001101";
		Trees_din <= x"030b980c";
		wait for Clk_period;
		Addr <=  "00000000001110";
		Trees_din <= x"03092d04";
		wait for Clk_period;
		Addr <=  "00000000001111";
		Trees_din <= x"ff540069";
		wait for Clk_period;
		Addr <=  "00000000010000";
		Trees_din <= x"00f0ae04";
		wait for Clk_period;
		Addr <=  "00000000010001";
		Trees_din <= x"ff620069";
		wait for Clk_period;
		Addr <=  "00000000010010";
		Trees_din <= x"01840069";
		wait for Clk_period;
		Addr <=  "00000000010011";
		Trees_din <= x"060d1808";
		wait for Clk_period;
		Addr <=  "00000000010100";
		Trees_din <= x"0609ea04";
		wait for Clk_period;
		Addr <=  "00000000010101";
		Trees_din <= x"01b90069";
		wait for Clk_period;
		Addr <=  "00000000010110";
		Trees_din <= x"00a60069";
		wait for Clk_period;
		Addr <=  "00000000010111";
		Trees_din <= x"0312d504";
		wait for Clk_period;
		Addr <=  "00000000011000";
		Trees_din <= x"ff610069";
		wait for Clk_period;
		Addr <=  "00000000011001";
		Trees_din <= x"01210069";
		wait for Clk_period;
		Addr <=  "00000000011010";
		Trees_din <= x"030b980c";
		wait for Clk_period;
		Addr <=  "00000000011011";
		Trees_din <= x"03092d04";
		wait for Clk_period;
		Addr <=  "00000000011100";
		Trees_din <= x"ff59009d";
		wait for Clk_period;
		Addr <=  "00000000011101";
		Trees_din <= x"00f0ae04";
		wait for Clk_period;
		Addr <=  "00000000011110";
		Trees_din <= x"ff68009d";
		wait for Clk_period;
		Addr <=  "00000000011111";
		Trees_din <= x"011d009d";
		wait for Clk_period;
		Addr <=  "00000000100000";
		Trees_din <= x"0613800c";
		wait for Clk_period;
		Addr <=  "00000000100001";
		Trees_din <= x"050e0408";
		wait for Clk_period;
		Addr <=  "00000000100010";
		Trees_din <= x"00c00004";
		wait for Clk_period;
		Addr <=  "00000000100011";
		Trees_din <= x"ffab009d";
		wait for Clk_period;
		Addr <=  "00000000100100";
		Trees_din <= x"013d009d";
		wait for Clk_period;
		Addr <=  "00000000100101";
		Trees_din <= x"ff92009d";
		wait for Clk_period;
		Addr <=  "00000000100110";
		Trees_din <= x"ff6b009d";
		wait for Clk_period;
		Addr <=  "00000000100111";
		Trees_din <= x"030b980c";
		wait for Clk_period;
		Addr <=  "00000000101000";
		Trees_din <= x"03092d04";
		wait for Clk_period;
		Addr <=  "00000000101001";
		Trees_din <= x"ff5c00d9";
		wait for Clk_period;
		Addr <=  "00000000101010";
		Trees_din <= x"00f0ae04";
		wait for Clk_period;
		Addr <=  "00000000101011";
		Trees_din <= x"ff6e00d9";
		wait for Clk_period;
		Addr <=  "00000000101100";
		Trees_din <= x"00e200d9";
		wait for Clk_period;
		Addr <=  "00000000101101";
		Trees_din <= x"06138010";
		wait for Clk_period;
		Addr <=  "00000000101110";
		Trees_din <= x"050e040c";
		wait for Clk_period;
		Addr <=  "00000000101111";
		Trees_din <= x"0100fc04";
		wait for Clk_period;
		Addr <=  "00000000110000";
		Trees_din <= x"010000d9";
		wait for Clk_period;
		Addr <=  "00000000110001";
		Trees_din <= x"09027404";
		wait for Clk_period;
		Addr <=  "00000000110010";
		Trees_din <= x"00a000d9";
		wait for Clk_period;
		Addr <=  "00000000110011";
		Trees_din <= x"fffe00d9";
		wait for Clk_period;
		Addr <=  "00000000110100";
		Trees_din <= x"ff9d00d9";
		wait for Clk_period;
		Addr <=  "00000000110101";
		Trees_din <= x"ff7200d9";
		wait for Clk_period;
		Addr <=  "00000000110110";
		Trees_din <= x"030b980c";
		wait for Clk_period;
		Addr <=  "00000000110111";
		Trees_din <= x"03092d04";
		wait for Clk_period;
		Addr <=  "00000000111000";
		Trees_din <= x"ff5f010d";
		wait for Clk_period;
		Addr <=  "00000000111001";
		Trees_din <= x"00f0ae04";
		wait for Clk_period;
		Addr <=  "00000000111010";
		Trees_din <= x"ff74010d";
		wait for Clk_period;
		Addr <=  "00000000111011";
		Trees_din <= x"00bc010d";
		wait for Clk_period;
		Addr <=  "00000000111100";
		Trees_din <= x"0613800c";
		wait for Clk_period;
		Addr <=  "00000000111101";
		Trees_din <= x"0100fc04";
		wait for Clk_period;
		Addr <=  "00000000111110";
		Trees_din <= x"00db010d";
		wait for Clk_period;
		Addr <=  "00000000111111";
		Trees_din <= x"060d1804";
		wait for Clk_period;
		Addr <=  "00000001000000";
		Trees_din <= x"007f010d";
		wait for Clk_period;
		Addr <=  "00000001000001";
		Trees_din <= x"ffa5010d";
		wait for Clk_period;
		Addr <=  "00000001000010";
		Trees_din <= x"ff78010d";
		wait for Clk_period;
		Addr <=  "00000001000011";
		Trees_din <= x"030b980c";
		wait for Clk_period;
		Addr <=  "00000001000100";
		Trees_din <= x"03092d04";
		wait for Clk_period;
		Addr <=  "00000001000101";
		Trees_din <= x"ff610141";
		wait for Clk_period;
		Addr <=  "00000001000110";
		Trees_din <= x"00f0ae04";
		wait for Clk_period;
		Addr <=  "00000001000111";
		Trees_din <= x"ff7b0141";
		wait for Clk_period;
		Addr <=  "00000001001000";
		Trees_din <= x"00a10141";
		wait for Clk_period;
		Addr <=  "00000001001001";
		Trees_din <= x"0613800c";
		wait for Clk_period;
		Addr <=  "00000001001010";
		Trees_din <= x"0100fc04";
		wait for Clk_period;
		Addr <=  "00000001001011";
		Trees_din <= x"00c50141";
		wait for Clk_period;
		Addr <=  "00000001001100";
		Trees_din <= x"0312d504";
		wait for Clk_period;
		Addr <=  "00000001001101";
		Trees_din <= x"ffd00141";
		wait for Clk_period;
		Addr <=  "00000001001110";
		Trees_din <= x"00820141";
		wait for Clk_period;
		Addr <=  "00000001001111";
		Trees_din <= x"ff7e0141";
		wait for Clk_period;
		Addr <=  "00000001010000";
		Trees_din <= x"030b980c";
		wait for Clk_period;
		Addr <=  "00000001010001";
		Trees_din <= x"03092d04";
		wait for Clk_period;
		Addr <=  "00000001010010";
		Trees_din <= x"ff630175";
		wait for Clk_period;
		Addr <=  "00000001010011";
		Trees_din <= x"00f0ae04";
		wait for Clk_period;
		Addr <=  "00000001010100";
		Trees_din <= x"ff820175";
		wait for Clk_period;
		Addr <=  "00000001010101";
		Trees_din <= x"008d0175";
		wait for Clk_period;
		Addr <=  "00000001010110";
		Trees_din <= x"040b520c";
		wait for Clk_period;
		Addr <=  "00000001010111";
		Trees_din <= x"0100fc04";
		wait for Clk_period;
		Addr <=  "00000001011000";
		Trees_din <= x"00b40175";
		wait for Clk_period;
		Addr <=  "00000001011001";
		Trees_din <= x"11024f04";
		wait for Clk_period;
		Addr <=  "00000001011010";
		Trees_din <= x"ffde0175";
		wait for Clk_period;
		Addr <=  "00000001011011";
		Trees_din <= x"00770175";
		wait for Clk_period;
		Addr <=  "00000001011100";
		Trees_din <= x"ff840175";
		wait for Clk_period;
		Addr <=  "00000001011101";
		Trees_din <= x"030b9814";
		wait for Clk_period;
		Addr <=  "00000001011110";
		Trees_din <= x"03092d0c";
		wait for Clk_period;
		Addr <=  "00000001011111";
		Trees_din <= x"03063404";
		wait for Clk_period;
		Addr <=  "00000001100000";
		Trees_din <= x"ff6301b9";
		wait for Clk_period;
		Addr <=  "00000001100001";
		Trees_din <= x"0605f104";
		wait for Clk_period;
		Addr <=  "00000001100010";
		Trees_din <= x"004601b9";
		wait for Clk_period;
		Addr <=  "00000001100011";
		Trees_din <= x"ff7d01b9";
		wait for Clk_period;
		Addr <=  "00000001100100";
		Trees_din <= x"00f0ae04";
		wait for Clk_period;
		Addr <=  "00000001100101";
		Trees_din <= x"ff8901b9";
		wait for Clk_period;
		Addr <=  "00000001100110";
		Trees_din <= x"007d01b9";
		wait for Clk_period;
		Addr <=  "00000001100111";
		Trees_din <= x"00c00004";
		wait for Clk_period;
		Addr <=  "00000001101000";
		Trees_din <= x"ff8a01b9";
		wait for Clk_period;
		Addr <=  "00000001101001";
		Trees_din <= x"0100fc04";
		wait for Clk_period;
		Addr <=  "00000001101010";
		Trees_din <= x"00a801b9";
		wait for Clk_period;
		Addr <=  "00000001101011";
		Trees_din <= x"0312d504";
		wait for Clk_period;
		Addr <=  "00000001101100";
		Trees_din <= x"ffe301b9";
		wait for Clk_period;
		Addr <=  "00000001101101";
		Trees_din <= x"006c01b9";
		wait for Clk_period;
		Addr <=  "00000001101110";
		Trees_din <= x"030b9810";
		wait for Clk_period;
		Addr <=  "00000001101111";
		Trees_din <= x"03063404";
		wait for Clk_period;
		Addr <=  "00000001110000";
		Trees_din <= x"ff6401f5";
		wait for Clk_period;
		Addr <=  "00000001110001";
		Trees_din <= x"00f6eb04";
		wait for Clk_period;
		Addr <=  "00000001110010";
		Trees_din <= x"ff7801f5";
		wait for Clk_period;
		Addr <=  "00000001110011";
		Trees_din <= x"13fafb04";
		wait for Clk_period;
		Addr <=  "00000001110100";
		Trees_din <= x"00ce01f5";
		wait for Clk_period;
		Addr <=  "00000001110101";
		Trees_din <= x"000d01f5";
		wait for Clk_period;
		Addr <=  "00000001110110";
		Trees_din <= x"0613800c";
		wait for Clk_period;
		Addr <=  "00000001110111";
		Trees_din <= x"0100fc04";
		wait for Clk_period;
		Addr <=  "00000001111000";
		Trees_din <= x"00a101f5";
		wait for Clk_period;
		Addr <=  "00000001111001";
		Trees_din <= x"05ff7004";
		wait for Clk_period;
		Addr <=  "00000001111010";
		Trees_din <= x"006201f5";
		wait for Clk_period;
		Addr <=  "00000001111011";
		Trees_din <= x"ffd601f5";
		wait for Clk_period;
		Addr <=  "00000001111100";
		Trees_din <= x"ff9101f5";
		wait for Clk_period;
		Addr <=  "00000001111101";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00000001111110";
		Trees_din <= x"030b980c";
		wait for Clk_period;
		Addr <=  "00000001111111";
		Trees_din <= x"03063404";
		wait for Clk_period;
		Addr <=  "00000010000000";
		Trees_din <= x"ff650225";
		wait for Clk_period;
		Addr <=  "00000010000001";
		Trees_din <= x"00f6eb04";
		wait for Clk_period;
		Addr <=  "00000010000010";
		Trees_din <= x"ff7d0225";
		wait for Clk_period;
		Addr <=  "00000010000011";
		Trees_din <= x"00870225";
		wait for Clk_period;
		Addr <=  "00000010000100";
		Trees_din <= x"040b5208";
		wait for Clk_period;
		Addr <=  "00000010000101";
		Trees_din <= x"05098d04";
		wait for Clk_period;
		Addr <=  "00000010000110";
		Trees_din <= x"00990225";
		wait for Clk_period;
		Addr <=  "00000010000111";
		Trees_din <= x"002a0225";
		wait for Clk_period;
		Addr <=  "00000010001000";
		Trees_din <= x"ff980225";
		wait for Clk_period;
		Addr <=  "00000010001001";
		Trees_din <= x"03092d0c";
		wait for Clk_period;
		Addr <=  "00000010001010";
		Trees_din <= x"03063404";
		wait for Clk_period;
		Addr <=  "00000010001011";
		Trees_din <= x"ff660259";
		wait for Clk_period;
		Addr <=  "00000010001100";
		Trees_din <= x"0b029504";
		wait for Clk_period;
		Addr <=  "00000010001101";
		Trees_din <= x"ff930259";
		wait for Clk_period;
		Addr <=  "00000010001110";
		Trees_din <= x"00480259";
		wait for Clk_period;
		Addr <=  "00000010001111";
		Trees_din <= x"0206390c";
		wait for Clk_period;
		Addr <=  "00000010010000";
		Trees_din <= x"0100fc08";
		wait for Clk_period;
		Addr <=  "00000010010001";
		Trees_din <= x"05098d04";
		wait for Clk_period;
		Addr <=  "00000010010010";
		Trees_din <= x"00990259";
		wait for Clk_period;
		Addr <=  "00000010010011";
		Trees_din <= x"00330259";
		wait for Clk_period;
		Addr <=  "00000010010100";
		Trees_din <= x"000a0259";
		wait for Clk_period;
		Addr <=  "00000010010101";
		Trees_din <= x"ff8d0259";
		wait for Clk_period;
		Addr <=  "00000010010110";
		Trees_din <= x"03092d0c";
		wait for Clk_period;
		Addr <=  "00000010010111";
		Trees_din <= x"03063404";
		wait for Clk_period;
		Addr <=  "00000010011000";
		Trees_din <= x"ff66028d";
		wait for Clk_period;
		Addr <=  "00000010011001";
		Trees_din <= x"02004104";
		wait for Clk_period;
		Addr <=  "00000010011010";
		Trees_din <= x"0047028d";
		wait for Clk_period;
		Addr <=  "00000010011011";
		Trees_din <= x"ff9b028d";
		wait for Clk_period;
		Addr <=  "00000010011100";
		Trees_din <= x"0206390c";
		wait for Clk_period;
		Addr <=  "00000010011101";
		Trees_din <= x"0100fc08";
		wait for Clk_period;
		Addr <=  "00000010011110";
		Trees_din <= x"05098d04";
		wait for Clk_period;
		Addr <=  "00000010011111";
		Trees_din <= x"0093028d";
		wait for Clk_period;
		Addr <=  "00000010100000";
		Trees_din <= x"002f028d";
		wait for Clk_period;
		Addr <=  "00000010100001";
		Trees_din <= x"000b028d";
		wait for Clk_period;
		Addr <=  "00000010100010";
		Trees_din <= x"ff95028d";
		wait for Clk_period;
		Addr <=  "00000010100011";
		Trees_din <= x"03063404";
		wait for Clk_period;
		Addr <=  "00000010100100";
		Trees_din <= x"ff6702b1";
		wait for Clk_period;
		Addr <=  "00000010100101";
		Trees_din <= x"0100fc08";
		wait for Clk_period;
		Addr <=  "00000010100110";
		Trees_din <= x"05098d04";
		wait for Clk_period;
		Addr <=  "00000010100111";
		Trees_din <= x"009002b1";
		wait for Clk_period;
		Addr <=  "00000010101000";
		Trees_din <= x"001a02b1";
		wait for Clk_period;
		Addr <=  "00000010101001";
		Trees_din <= x"060d1804";
		wait for Clk_period;
		Addr <=  "00000010101010";
		Trees_din <= x"000e02b1";
		wait for Clk_period;
		Addr <=  "00000010101011";
		Trees_din <= x"ff8902b1";
		wait for Clk_period;
		Addr <=  "00000010101100";
		Trees_din <= x"03063404";
		wait for Clk_period;
		Addr <=  "00000010101101";
		Trees_din <= x"ff6802d5";
		wait for Clk_period;
		Addr <=  "00000010101110";
		Trees_din <= x"0100fc08";
		wait for Clk_period;
		Addr <=  "00000010101111";
		Trees_din <= x"02ff7004";
		wait for Clk_period;
		Addr <=  "00000010110000";
		Trees_din <= x"008d02d5";
		wait for Clk_period;
		Addr <=  "00000010110001";
		Trees_din <= x"002302d5";
		wait for Clk_period;
		Addr <=  "00000010110010";
		Trees_din <= x"060d1804";
		wait for Clk_period;
		Addr <=  "00000010110011";
		Trees_din <= x"000d02d5";
		wait for Clk_period;
		Addr <=  "00000010110100";
		Trees_din <= x"ff9002d5";
		wait for Clk_period;
		Addr <=  "00000010110101";
		Trees_din <= x"03063404";
		wait for Clk_period;
		Addr <=  "00000010110110";
		Trees_din <= x"ff690301";
		wait for Clk_period;
		Addr <=  "00000010110111";
		Trees_din <= x"0100fc0c";
		wait for Clk_period;
		Addr <=  "00000010111000";
		Trees_din <= x"05098d08";
		wait for Clk_period;
		Addr <=  "00000010111001";
		Trees_din <= x"05fb3c04";
		wait for Clk_period;
		Addr <=  "00000010111010";
		Trees_din <= x"001f0301";
		wait for Clk_period;
		Addr <=  "00000010111011";
		Trees_din <= x"008c0301";
		wait for Clk_period;
		Addr <=  "00000010111100";
		Trees_din <= x"00110301";
		wait for Clk_period;
		Addr <=  "00000010111101";
		Trees_din <= x"04093c04";
		wait for Clk_period;
		Addr <=  "00000010111110";
		Trees_din <= x"000d0301";
		wait for Clk_period;
		Addr <=  "00000010111111";
		Trees_din <= x"ff980301";
		wait for Clk_period;
		Addr <=  "00000011000000";
		Trees_din <= x"03063404";
		wait for Clk_period;
		Addr <=  "00000011000001";
		Trees_din <= x"ff6a032d";
		wait for Clk_period;
		Addr <=  "00000011000010";
		Trees_din <= x"0609ea0c";
		wait for Clk_period;
		Addr <=  "00000011000011";
		Trees_din <= x"00e9ab04";
		wait for Clk_period;
		Addr <=  "00000011000100";
		Trees_din <= x"001a032d";
		wait for Clk_period;
		Addr <=  "00000011000101";
		Trees_din <= x"0d009204";
		wait for Clk_period;
		Addr <=  "00000011000110";
		Trees_din <= x"0025032d";
		wait for Clk_period;
		Addr <=  "00000011000111";
		Trees_din <= x"008a032d";
		wait for Clk_period;
		Addr <=  "00000011001000";
		Trees_din <= x"17004704";
		wait for Clk_period;
		Addr <=  "00000011001001";
		Trees_din <= x"ff9f032d";
		wait for Clk_period;
		Addr <=  "00000011001010";
		Trees_din <= x"0013032d";
		wait for Clk_period;
		Addr <=  "00000011001011";
		Trees_din <= x"03063404";
		wait for Clk_period;
		Addr <=  "00000011001100";
		Trees_din <= x"ff6b0351";
		wait for Clk_period;
		Addr <=  "00000011001101";
		Trees_din <= x"0206390c";
		wait for Clk_period;
		Addr <=  "00000011001110";
		Trees_din <= x"1e006504";
		wait for Clk_period;
		Addr <=  "00000011001111";
		Trees_din <= x"000b0351";
		wait for Clk_period;
		Addr <=  "00000011010000";
		Trees_din <= x"1e007704";
		wait for Clk_period;
		Addr <=  "00000011010001";
		Trees_din <= x"00840351";
		wait for Clk_period;
		Addr <=  "00000011010010";
		Trees_din <= x"00200351";
		wait for Clk_period;
		Addr <=  "00000011010011";
		Trees_din <= x"ffa50351";
		wait for Clk_period;
		Addr <=  "00000011010100";
		Trees_din <= x"03063404";
		wait for Clk_period;
		Addr <=  "00000011010101";
		Trees_din <= x"ff6d0375";
		wait for Clk_period;
		Addr <=  "00000011010110";
		Trees_din <= x"0100fc08";
		wait for Clk_period;
		Addr <=  "00000011010111";
		Trees_din <= x"02fe0004";
		wait for Clk_period;
		Addr <=  "00000011011000";
		Trees_din <= x"00700375";
		wait for Clk_period;
		Addr <=  "00000011011001";
		Trees_din <= x"00100375";
		wait for Clk_period;
		Addr <=  "00000011011010";
		Trees_din <= x"00c00004";
		wait for Clk_period;
		Addr <=  "00000011011011";
		Trees_din <= x"ffae0375";
		wait for Clk_period;
		Addr <=  "00000011011100";
		Trees_din <= x"fffc0375";
		wait for Clk_period;
		Addr <=  "00000011011101";
		Trees_din <= x"03063404";
		wait for Clk_period;
		Addr <=  "00000011011110";
		Trees_din <= x"ff6f0391";
		wait for Clk_period;
		Addr <=  "00000011011111";
		Trees_din <= x"040b5208";
		wait for Clk_period;
		Addr <=  "00000011100000";
		Trees_din <= x"030d7004";
		wait for Clk_period;
		Addr <=  "00000011100001";
		Trees_din <= x"000c0391";
		wait for Clk_period;
		Addr <=  "00000011100010";
		Trees_din <= x"00660391";
		wait for Clk_period;
		Addr <=  "00000011100011";
		Trees_din <= x"ffb10391";
		wait for Clk_period;
		Addr <=  "00000011100100";
		Trees_din <= x"03063404";
		wait for Clk_period;
		Addr <=  "00000011100101";
		Trees_din <= x"ff7103ad";
		wait for Clk_period;
		Addr <=  "00000011100110";
		Trees_din <= x"0100fc08";
		wait for Clk_period;
		Addr <=  "00000011100111";
		Trees_din <= x"02fe0004";
		wait for Clk_period;
		Addr <=  "00000011101000";
		Trees_din <= x"006103ad";
		wait for Clk_period;
		Addr <=  "00000011101001";
		Trees_din <= x"000703ad";
		wait for Clk_period;
		Addr <=  "00000011101010";
		Trees_din <= x"ffce03ad";
		wait for Clk_period;
		Addr <=  "00000011101011";
		Trees_din <= x"03063404";
		wait for Clk_period;
		Addr <=  "00000011101100";
		Trees_din <= x"ff7403c9";
		wait for Clk_period;
		Addr <=  "00000011101101";
		Trees_din <= x"0609ea08";
		wait for Clk_period;
		Addr <=  "00000011101110";
		Trees_din <= x"06fed504";
		wait for Clk_period;
		Addr <=  "00000011101111";
		Trees_din <= x"000c03c9";
		wait for Clk_period;
		Addr <=  "00000011110000";
		Trees_din <= x"005f03c9";
		wait for Clk_period;
		Addr <=  "00000011110001";
		Trees_din <= x"ffd803c9";
		wait for Clk_period;
		Addr <=  "00000011110010";
		Trees_din <= x"03063404";
		wait for Clk_period;
		Addr <=  "00000011110011";
		Trees_din <= x"ff7703e5";
		wait for Clk_period;
		Addr <=  "00000011110100";
		Trees_din <= x"02ff7008";
		wait for Clk_period;
		Addr <=  "00000011110101";
		Trees_din <= x"08005504";
		wait for Clk_period;
		Addr <=  "00000011110110";
		Trees_din <= x"001203e5";
		wait for Clk_period;
		Addr <=  "00000011110111";
		Trees_din <= x"005b03e5";
		wait for Clk_period;
		Addr <=  "00000011111000";
		Trees_din <= x"ffdc03e5";
		wait for Clk_period;
		Addr <=  "00000011111001";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00000011111010";
		Trees_din <= x"03063404";
		wait for Clk_period;
		Addr <=  "00000011111011";
		Trees_din <= x"ff7a0405";
		wait for Clk_period;
		Addr <=  "00000011111100";
		Trees_din <= x"0312d508";
		wait for Clk_period;
		Addr <=  "00000011111101";
		Trees_din <= x"00e9ab04";
		wait for Clk_period;
		Addr <=  "00000011111110";
		Trees_din <= x"ffab0405";
		wait for Clk_period;
		Addr <=  "00000011111111";
		Trees_din <= x"00370405";
		wait for Clk_period;
		Addr <=  "00000100000000";
		Trees_din <= x"00580405";
		wait for Clk_period;
		Addr <=  "00000100000001";
		Trees_din <= x"030d7008";
		wait for Clk_period;
		Addr <=  "00000100000010";
		Trees_din <= x"07004f04";
		wait for Clk_period;
		Addr <=  "00000100000011";
		Trees_din <= x"fffd0419";
		wait for Clk_period;
		Addr <=  "00000100000100";
		Trees_din <= x"ff830419";
		wait for Clk_period;
		Addr <=  "00000100000101";
		Trees_din <= x"00460419";
		wait for Clk_period;
		Addr <=  "00000100000110";
		Trees_din <= x"03063404";
		wait for Clk_period;
		Addr <=  "00000100000111";
		Trees_din <= x"ff82042d";
		wait for Clk_period;
		Addr <=  "00000100001000";
		Trees_din <= x"02ff7004";
		wait for Clk_period;
		Addr <=  "00000100001001";
		Trees_din <= x"0040042d";
		wait for Clk_period;
		Addr <=  "00000100001010";
		Trees_din <= x"ffe6042d";
		wait for Clk_period;
		Addr <=  "00000100001011";
		Trees_din <= x"03063404";
		wait for Clk_period;
		Addr <=  "00000100001100";
		Trees_din <= x"ff870441";
		wait for Clk_period;
		Addr <=  "00000100001101";
		Trees_din <= x"02ff7004";
		wait for Clk_period;
		Addr <=  "00000100001110";
		Trees_din <= x"003a0441";
		wait for Clk_period;
		Addr <=  "00000100001111";
		Trees_din <= x"ffe80441";
		wait for Clk_period;
		Addr <=  "00000100010000";
		Trees_din <= x"030d7008";
		wait for Clk_period;
		Addr <=  "00000100010001";
		Trees_din <= x"03063404";
		wait for Clk_period;
		Addr <=  "00000100010010";
		Trees_din <= x"ff8c0455";
		wait for Clk_period;
		Addr <=  "00000100010011";
		Trees_din <= x"ffec0455";
		wait for Clk_period;
		Addr <=  "00000100010100";
		Trees_din <= x"003d0455";
		wait for Clk_period;
		Addr <=  "00000100010101";
		Trees_din <= x"030d7008";
		wait for Clk_period;
		Addr <=  "00000100010110";
		Trees_din <= x"03063404";
		wait for Clk_period;
		Addr <=  "00000100010111";
		Trees_din <= x"ff910469";
		wait for Clk_period;
		Addr <=  "00000100011000";
		Trees_din <= x"ffee0469";
		wait for Clk_period;
		Addr <=  "00000100011001";
		Trees_din <= x"00380469";
		wait for Clk_period;
		Addr <=  "00000100011010";
		Trees_din <= x"030d7008";
		wait for Clk_period;
		Addr <=  "00000100011011";
		Trees_din <= x"03063404";
		wait for Clk_period;
		Addr <=  "00000100011100";
		Trees_din <= x"ff96047d";
		wait for Clk_period;
		Addr <=  "00000100011101";
		Trees_din <= x"ffef047d";
		wait for Clk_period;
		Addr <=  "00000100011110";
		Trees_din <= x"0034047d";
		wait for Clk_period;
		Addr <=  "00000100011111";
		Trees_din <= x"030b9808";
		wait for Clk_period;
		Addr <=  "00000100100000";
		Trees_din <= x"15fa8d04";
		wait for Clk_period;
		Addr <=  "00000100100001";
		Trees_din <= x"ffec0491";
		wait for Clk_period;
		Addr <=  "00000100100010";
		Trees_din <= x"ff9e0491";
		wait for Clk_period;
		Addr <=  "00000100100011";
		Trees_din <= x"002b0491";
		wait for Clk_period;
		Addr <=  "00000100100100";
		Trees_din <= x"03063404";
		wait for Clk_period;
		Addr <=  "00000100100101";
		Trees_din <= x"ff9f04a5";
		wait for Clk_period;
		Addr <=  "00000100100110";
		Trees_din <= x"02fbc304";
		wait for Clk_period;
		Addr <=  "00000100100111";
		Trees_din <= x"003104a5";
		wait for Clk_period;
		Addr <=  "00000100101000";
		Trees_din <= x"ffef04a5";
		wait for Clk_period;
		Addr <=  "00000100101001";
		Trees_din <= x"03017804";
		wait for Clk_period;
		Addr <=  "00000100101010";
		Trees_din <= x"ffa804b9";
		wait for Clk_period;
		Addr <=  "00000100101011";
		Trees_din <= x"12009204";
		wait for Clk_period;
		Addr <=  "00000100101100";
		Trees_din <= x"002604b9";
		wait for Clk_period;
		Addr <=  "00000100101101";
		Trees_din <= x"ffea04b9";
		wait for Clk_period;
		Addr <=  "00000100101110";
		Trees_din <= x"03017804";
		wait for Clk_period;
		Addr <=  "00000100101111";
		Trees_din <= x"ffad04cd";
		wait for Clk_period;
		Addr <=  "00000100110000";
		Trees_din <= x"13fb5504";
		wait for Clk_period;
		Addr <=  "00000100110001";
		Trees_din <= x"002004cd";
		wait for Clk_period;
		Addr <=  "00000100110010";
		Trees_din <= x"fff004cd";
		wait for Clk_period;
		Addr <=  "00000100110011";
		Trees_din <= x"02fbc304";
		wait for Clk_period;
		Addr <=  "00000100110100";
		Trees_din <= x"001a04d9";
		wait for Clk_period;
		Addr <=  "00000100110101";
		Trees_din <= x"ffc104d9";
		wait for Clk_period;
		Addr <=  "00000100110110";
		Trees_din <= x"030b9804";
		wait for Clk_period;
		Addr <=  "00000100110111";
		Trees_din <= x"ffbb04e5";
		wait for Clk_period;
		Addr <=  "00000100111000";
		Trees_din <= x"002804e5";
		wait for Clk_period;
		Addr <=  "00000100111001";
		Trees_din <= x"02fcdf04";
		wait for Clk_period;
		Addr <=  "00000100111010";
		Trees_din <= x"001504f1";
		wait for Clk_period;
		Addr <=  "00000100111011";
		Trees_din <= x"ffcb04f1";
		wait for Clk_period;
		Addr <=  "00000100111100";
		Trees_din <= x"03092d04";
		wait for Clk_period;
		Addr <=  "00000100111101";
		Trees_din <= x"ffbf04fd";
		wait for Clk_period;
		Addr <=  "00000100111110";
		Trees_din <= x"002504fd";
		wait for Clk_period;
		Addr <=  "00000100111111";
		Trees_din <= x"02fe0004";
		wait for Clk_period;
		Addr <=  "00000101000000";
		Trees_din <= x"00120509";
		wait for Clk_period;
		Addr <=  "00000101000001";
		Trees_din <= x"ffce0509";
		wait for Clk_period;
		Addr <=  "00000101000010";
		Trees_din <= x"02fe0004";
		wait for Clk_period;
		Addr <=  "00000101000011";
		Trees_din <= x"00110515";
		wait for Clk_period;
		Addr <=  "00000101000100";
		Trees_din <= x"ffd10515";
		wait for Clk_period;
		Addr <=  "00000101000101";
		Trees_din <= x"02fe0004";
		wait for Clk_period;
		Addr <=  "00000101000110";
		Trees_din <= x"00100521";
		wait for Clk_period;
		Addr <=  "00000101000111";
		Trees_din <= x"ffd40521";
		wait for Clk_period;
		Addr <=  "00000101001000";
		Trees_din <= x"12009304";
		wait for Clk_period;
		Addr <=  "00000101001001";
		Trees_din <= x"000d052d";
		wait for Clk_period;
		Addr <=  "00000101001010";
		Trees_din <= x"ffd8052d";
		wait for Clk_period;
		Addr <=  "00000101001011";
		Trees_din <= x"17004504";
		wait for Clk_period;
		Addr <=  "00000101001100";
		Trees_din <= x"ffdb0539";
		wait for Clk_period;
		Addr <=  "00000101001101";
		Trees_din <= x"000c0539";
		wait for Clk_period;
		Addr <=  "00000101001110";
		Trees_din <= x"0b013604";
		wait for Clk_period;
		Addr <=  "00000101001111";
		Trees_din <= x"ffe60545";
		wait for Clk_period;
		Addr <=  "00000101010000";
		Trees_din <= x"00030545";
		wait for Clk_period;
		Addr <=  "00000101010001";
		Trees_din <= x"fff20549";
		wait for Clk_period;
		Addr <=  "00000101010010";
		Trees_din <= x"fff2054d";
		wait for Clk_period;
		Addr <=  "00000101010011";
		Trees_din <= x"fff40551";
		wait for Clk_period;
		Addr <=  "00000101010100";
		Trees_din <= x"fff40555";
		wait for Clk_period;
		Addr <=  "00000101010101";
		Trees_din <= x"fff60559";
		wait for Clk_period;
		Addr <=  "00000101010110";
		Trees_din <= x"fff6055d";
		wait for Clk_period;
		Addr <=  "00000101010111";
		Trees_din <= x"fff70561";
		wait for Clk_period;
		Addr <=  "00000101011000";
		Trees_din <= x"fff70565";
		wait for Clk_period;
		Addr <=  "00000101011001";
		Trees_din <= x"fff80569";
		wait for Clk_period;
		Addr <=  "00000101011010";
		Trees_din <= x"fff9056d";
		wait for Clk_period;
		Addr <=  "00000101011011";
		Trees_din <= x"fff90571";
		wait for Clk_period;
		Addr <=  "00000101011100";
		Trees_din <= x"fff90575";
		wait for Clk_period;
		Addr <=  "00000101011101";
		Trees_din <= x"fff90579";
		wait for Clk_period;
		Addr <=  "00000101011110";
		Trees_din <= x"fffa057d";
		wait for Clk_period;
		Addr <=  "00000101011111";
		Trees_din <= x"fffa0581";
		wait for Clk_period;
		Addr <=  "00000101100000";
		Trees_din <= x"fffa0585";
		wait for Clk_period;
		Addr <=  "00000101100001";
		Trees_din <= x"fffb0589";
		wait for Clk_period;
		Addr <=  "00000101100010";
		Trees_din <= x"fffc058d";
		wait for Clk_period;
		Addr <=  "00000101100011";
		Trees_din <= x"fffb0591";
		wait for Clk_period;
		Addr <=  "00000101100100";
		Trees_din <= x"fffb0595";
		wait for Clk_period;
		Addr <=  "00000101100101";
		Trees_din <= x"fffb0599";
		wait for Clk_period;
		Addr <=  "00000101100110";
		Trees_din <= x"fffc059d";
		wait for Clk_period;
		Addr <=  "00000101100111";
		Trees_din <= x"fffc05a1";
		wait for Clk_period;
		Addr <=  "00000101101000";
		Trees_din <= x"fffc05a5";
		wait for Clk_period;
		Addr <=  "00000101101001";
		Trees_din <= x"fffc05a9";
		wait for Clk_period;
		Addr <=  "00000101101010";
		Trees_din <= x"fffd05ad";
		wait for Clk_period;
		Addr <=  "00000101101011";
		Trees_din <= x"fffc05b1";
		wait for Clk_period;
		Addr <=  "00000101101100";
		Trees_din <= x"fffc05b5";
		wait for Clk_period;
		Addr <=  "00000101101101";
		Trees_din <= x"fffd05b9";
		wait for Clk_period;
		Addr <=  "00000101101110";
		Trees_din <= x"fffd05bd";
		wait for Clk_period;
		Addr <=  "00000101101111";
		Trees_din <= x"fffd05c1";
		wait for Clk_period;
		Addr <=  "00000101110000";
		Trees_din <= x"fffd05c5";
		wait for Clk_period;
		Addr <=  "00000101110001";
		Trees_din <= x"fffe05c9";
		wait for Clk_period;
		Addr <=  "00000101110010";
		Trees_din <= x"fffe05cd";
		wait for Clk_period;
		Addr <=  "00000101110011";
		Trees_din <= x"fffe05d1";
		wait for Clk_period;
		Addr <=  "00000101110100";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00000101110101";
		Trees_din <= x"fffe05d9";
		wait for Clk_period;
		Addr <=  "00000101110110";
		Trees_din <= x"0000001f";
		wait for Clk_period;

        -- Reset valid flag
        Valid_node <= '0';
        wait for Clk_period; 
        
        class_label <= std_logic_vector(to_unsigned(5, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110101100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "0000001010010111";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "0000001011111110";
        wait for Clk_period; 
        Features_din <= "0000001000001100";
        wait for Clk_period; 
        Features_din <= "0000000111001000";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000010100011100";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000001000101101";
        wait for Clk_period; 
        Features_din <= "0000000100111011";
        wait for Clk_period; 
        Features_din <= "0000000011011110";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "0000001010100110";
        wait for Clk_period; 
        Features_din <= "0000001000001101";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "1111101100000001";
        wait for Clk_period; 
        Features_din <= "0000001100010101";
        wait for Clk_period; 
        Features_din <= "1111100101001101";
        wait for Clk_period; 
        Features_din <= "0000000100010010";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110110101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "0000001001110110";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000001100010110";
        wait for Clk_period; 
        Features_din <= "0000001001000001";
        wait for Clk_period; 
        Features_din <= "0000001000001001";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000001010001000";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111100110100101";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "1111100110110101";
        wait for Clk_period; 
        Features_din <= "0000001010001000";
        wait for Clk_period; 
        Features_din <= "0000001010001000";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "0000001010001000";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001010001000";
        wait for Clk_period; 
        Features_din <= "0000000011111100";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000110001110";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001010110101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "0000001000111100";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "0000001011001011";
        wait for Clk_period; 
        Features_din <= "0000001000101001";
        wait for Clk_period; 
        Features_din <= "0000000110010011";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111100010000111";
        wait for Clk_period; 
        Features_din <= "0000000011101101";
        wait for Clk_period; 
        Features_din <= "0000010100100111";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000000011100110";
        wait for Clk_period; 
        Features_din <= "1111110101011001";
        wait for Clk_period; 
        Features_din <= "0000000110101011";
        wait for Clk_period; 
        Features_din <= "1111111001010111";
        wait for Clk_period; 
        Features_din <= "0000000100100101";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000000011110010";
        wait for Clk_period; 
        Features_din <= "0000000110110011";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000001000100111";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000011101001";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111110000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011001100";
        wait for Clk_period; 
        Features_din <= "0000001001010110";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "0000001100011001";
        wait for Clk_period; 
        Features_din <= "0000001000000101";
        wait for Clk_period; 
        Features_din <= "0000000111110001";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000010010100111";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "1111111001000011";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "1111100011010000";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111000000011";
        wait for Clk_period; 
        Features_din <= "0000001010111010";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "0000000111111100";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010100110001";
        wait for Clk_period; 
        Features_din <= "0000001011010011";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110011010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "0000001001011011";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001001000111";
        wait for Clk_period; 
        Features_din <= "0000000111110011";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "1111011011111011";
        wait for Clk_period; 
        Features_din <= "0000000101011100";
        wait for Clk_period; 
        Features_din <= "0000000100001000";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "0000000110001010";
        wait for Clk_period; 
        Features_din <= "0000000100011001";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000000110110011";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001000010111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011101000";
        wait for Clk_period; 
        Features_din <= "0000001001000110";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001000001110";
        wait for Clk_period; 
        Features_din <= "0000000111110011";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000010100000000";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "1111111001001010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "1111100010100000";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111110111110101";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000111001000";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000011000000";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001001010010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "0000001000110111";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "0000001011111001";
        wait for Clk_period; 
        Features_din <= "0000001000110100";
        wait for Clk_period; 
        Features_din <= "0000000111010001";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000010100100011";
        wait for Clk_period; 
        Features_din <= "0000001000110010";
        wait for Clk_period; 
        Features_din <= "1111110100011110";
        wait for Clk_period; 
        Features_din <= "0000000100001010";
        wait for Clk_period; 
        Features_din <= "0000000111011111";
        wait for Clk_period; 
        Features_din <= "1111100101000110";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111001100110";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "0000000100110001";
        wait for Clk_period; 
        Features_din <= "0000000101010110";
        wait for Clk_period; 
        Features_din <= "0000010101001001";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000001100010001";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000011100101";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110001011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "0000001000110011";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001000101010";
        wait for Clk_period; 
        Features_din <= "0000000111100110";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000010010000110";
        wait for Clk_period; 
        Features_din <= "0000001000011100";
        wait for Clk_period; 
        Features_din <= "0000011001000111";
        wait for Clk_period; 
        Features_din <= "0000000111011011";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "1111110011001111";
        wait for Clk_period; 
        Features_din <= "0000000101000011";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "0000000100101000";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "1111101010110001";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "1111110010000011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000010111111";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111001100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "0000001001011000";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "0000001011100001";
        wait for Clk_period; 
        Features_din <= "0000001001100100";
        wait for Clk_period; 
        Features_din <= "0000001000000000";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "1111100111110011";
        wait for Clk_period; 
        Features_din <= "0000000101111100";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "1111100101101001";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000011001000";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000011011101";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110100011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "0000001001101011";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "0000001100110001";
        wait for Clk_period; 
        Features_din <= "0000001000100110";
        wait for Clk_period; 
        Features_din <= "0000001000001011";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000010011111010";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000001001110100";
        wait for Clk_period; 
        Features_din <= "0000000101111100";
        wait for Clk_period; 
        Features_din <= "1111110101000100";
        wait for Clk_period; 
        Features_din <= "0000000111010100";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "0000000101111111";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "1111100000010001";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001001011011";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000001000100010";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000011001011";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111010101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "0000001001011001";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000001100101000";
        wait for Clk_period; 
        Features_din <= "0000000111110001";
        wait for Clk_period; 
        Features_din <= "0000000111110010";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111111000000111";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111100000001110";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "0000000011001001";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111010100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "0000001001010110";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000001100001011";
        wait for Clk_period; 
        Features_din <= "0000001000011010";
        wait for Clk_period; 
        Features_din <= "0000000111011101";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111101000001000";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000000101000100";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000011000100001";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000000100111110";
        wait for Clk_period; 
        Features_din <= "0000000011010101";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111101101100010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000001001011001";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000011001000";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111111000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "0000001100110010";
        wait for Clk_period; 
        Features_din <= "0000001001011100";
        wait for Clk_period; 
        Features_din <= "0000000111011100";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "1111011101000001";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000001001110000";
        wait for Clk_period; 
        Features_din <= "1111111000111110";
        wait for Clk_period; 
        Features_din <= "0000000101111000";
        wait for Clk_period; 
        Features_din <= "0000000100101000";
        wait for Clk_period; 
        Features_din <= "0000001100101001";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000001010010000";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000010010110000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000011100110";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010111100";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001000101010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "0000001001011011";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000001100001101";
        wait for Clk_period; 
        Features_din <= "0000001000011001";
        wait for Clk_period; 
        Features_din <= "0000000111110001";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111100101011000";
        wait for Clk_period; 
        Features_din <= "0000000100001001";
        wait for Clk_period; 
        Features_din <= "0000000111010111";
        wait for Clk_period; 
        Features_din <= "0000000011111000";
        wait for Clk_period; 
        Features_din <= "0000000100000111";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "0000001010000000";
        wait for Clk_period; 
        Features_din <= "0000001000100100";
        wait for Clk_period; 
        Features_din <= "0000001010010010";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "1111101100001100";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010101011111";
        wait for Clk_period; 
        Features_din <= "0000001010111000";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000110111000";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111100110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010111101";
        wait for Clk_period; 
        Features_din <= "0000001000110101";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "0000001100101001";
        wait for Clk_period; 
        Features_din <= "0000001000011000";
        wait for Clk_period; 
        Features_din <= "0000000111010110";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "1111101010110100";
        wait for Clk_period; 
        Features_din <= "0000000011001000";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000000010101100";
        wait for Clk_period; 
        Features_din <= "0000000100111000";
        wait for Clk_period; 
        Features_din <= "0000000110001001";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "1111110011001111";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "1111101100010110";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000111001001";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001000111001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "0000001001011111";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000001100001110";
        wait for Clk_period; 
        Features_din <= "0000001000000100";
        wait for Clk_period; 
        Features_din <= "0000000111000101";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000010100100100";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111110110100110";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111100100011000";
        wait for Clk_period; 
        Features_din <= "1111111010101000";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "0000001010110000";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000110010110";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010100100100";
        wait for Clk_period; 
        Features_din <= "0000001011110100";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000100011100";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110110011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010111001";
        wait for Clk_period; 
        Features_din <= "0000001000110000";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001000111011";
        wait for Clk_period; 
        Features_din <= "0000001000011001";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001011101101";
        wait for Clk_period; 
        Features_din <= "1111100110000011";
        wait for Clk_period; 
        Features_din <= "0000001001101011";
        wait for Clk_period; 
        Features_din <= "0000001011000011";
        wait for Clk_period; 
        Features_din <= "1111100111010111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000000110010111";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001000000011";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000111011000";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000011100110";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111001101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "0000001001011111";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000001000011011";
        wait for Clk_period; 
        Features_din <= "0000000111110010";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111110110100000";
        wait for Clk_period; 
        Features_din <= "0000000101001110";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "0000000111010000";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000000101100100";
        wait for Clk_period; 
        Features_din <= "1111101101101101";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001010100110";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "1111101101111110";
        wait for Clk_period; 
        Features_din <= "0000001100000110";
        wait for Clk_period; 
        Features_din <= "0000011100010001";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000001001000101";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111100101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "0000001001010010";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000001100100010";
        wait for Clk_period; 
        Features_din <= "0000001000001001";
        wait for Clk_period; 
        Features_din <= "0000000111101101";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111110110101011";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111011111101110";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001000000100";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000011110011";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000011000100";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000101111111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "0000001001010000";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001000011010";
        wait for Clk_period; 
        Features_din <= "0000001000000100";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111100111011000";
        wait for Clk_period; 
        Features_din <= "0000000100010111";
        wait for Clk_period; 
        Features_din <= "0000001000110101";
        wait for Clk_period; 
        Features_din <= "0000000101111110";
        wait for Clk_period; 
        Features_din <= "0000001000101100";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000001001011100";
        wait for Clk_period; 
        Features_din <= "0000001100001101";
        wait for Clk_period; 
        Features_din <= "0000001011111010";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000000100111101";
        wait for Clk_period; 
        Features_din <= "1111100111111000";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000010101101";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000011100000";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111111101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "0000001001000111";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000001000000010";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000011001101011";
        wait for Clk_period; 
        Features_din <= "0000000100111011";
        wait for Clk_period; 
        Features_din <= "0000000111001111";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000001000111000";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "0000001000101010";
        wait for Clk_period; 
        Features_din <= "0000000101000010";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "1111101100101111";
        wait for Clk_period; 
        Features_din <= "0000001001001000";
        wait for Clk_period; 
        Features_din <= "1111100111011110";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000001100001100";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000010111111";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111101010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "0000001001001100";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000000111111001";
        wait for Clk_period; 
        Features_din <= "0000001000010011";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000011000000001";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "1111110110001011";
        wait for Clk_period; 
        Features_din <= "0000001100110011";
        wait for Clk_period; 
        Features_din <= "0000000111100101";
        wait for Clk_period; 
        Features_din <= "1111101110000101";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111110011111011";
        wait for Clk_period; 
        Features_din <= "0000000101011011";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "0000011000101111";
        wait for Clk_period; 
        Features_din <= "0000001001000011";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000001000111100";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110001100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "0000001001111001";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001000011100";
        wait for Clk_period; 
        Features_din <= "0000001000001000";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "1111110110011010";
        wait for Clk_period; 
        Features_din <= "0000000100101010";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000111001111";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111011111011100";
        wait for Clk_period; 
        Features_din <= "0000001011101010";
        wait for Clk_period; 
        Features_din <= "0000010011111100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000001010101111";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110001101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011100010";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001000100011";
        wait for Clk_period; 
        Features_din <= "0000001000010010";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000010011000100";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000011011001";
        wait for Clk_period; 
        Features_din <= "1111110111100110";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000011011010";
        wait for Clk_period; 
        Features_din <= "0000001011110011";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "1111011111010111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001001111101";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000110100000";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000000011010111";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111100001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "0000001000011100";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "0000001011110111";
        wait for Clk_period; 
        Features_din <= "0000001001001001";
        wait for Clk_period; 
        Features_din <= "0000000111011011";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "1111100111101101";
        wait for Clk_period; 
        Features_din <= "0000000100011011";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "1111100101101111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000011100110";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111100110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "0000001001111001";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "0000001100011110";
        wait for Clk_period; 
        Features_din <= "0000001000101011";
        wait for Clk_period; 
        Features_din <= "0000000111011111";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000001001000010";
        wait for Clk_period; 
        Features_din <= "0000001011101100";
        wait for Clk_period; 
        Features_din <= "0000000110011101";
        wait for Clk_period; 
        Features_din <= "0000000101110100";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000000011101011";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "1111101100100010";
        wait for Clk_period; 
        Features_din <= "0000000110000011";
        wait for Clk_period; 
        Features_din <= "1111100101101110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000001011101111";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000011011100";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110011101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "0000001100000100";
        wait for Clk_period; 
        Features_din <= "0000001000110000";
        wait for Clk_period; 
        Features_din <= "0000000111111011";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000111001011";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "1111111000001100";
        wait for Clk_period; 
        Features_din <= "0000000011110010";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "0000001000111011";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000001011110100";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "1111011101000001";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(3, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110001100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "0000001001100000";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000001100110001";
        wait for Clk_period; 
        Features_din <= "0000001000101111";
        wait for Clk_period; 
        Features_din <= "0000000111100010";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000101110111";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "1111110111010000";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "1111011110001010";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000000111011100";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000011110111";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000011010110";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001010000000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "0000001000111011";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "0000001011001010";
        wait for Clk_period; 
        Features_din <= "0000001000111001";
        wait for Clk_period; 
        Features_din <= "0000000111000111";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111101011100001";
        wait for Clk_period; 
        Features_din <= "0000000111011010";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000011100100";
        wait for Clk_period; 
        Features_din <= "0000000101011001";
        wait for Clk_period; 
        Features_din <= "0000010010010101";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "1111110011000111";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "1111101011111111";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000010111100";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110100111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "0000001010001010";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000001001001000";
        wait for Clk_period; 
        Features_din <= "0000001000000111";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "1111110100001001";
        wait for Clk_period; 
        Features_din <= "0000000101000000";
        wait for Clk_period; 
        Features_din <= "0000010101011111";
        wait for Clk_period; 
        Features_din <= "0000001000101011";
        wait for Clk_period; 
        Features_din <= "0000000101100000";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "0000010100111111";
        wait for Clk_period; 
        Features_din <= "0000000110011110";
        wait for Clk_period; 
        Features_din <= "0000001100010001";
        wait for Clk_period; 
        Features_din <= "0000000010101101";
        wait for Clk_period; 
        Features_din <= "1111110000101101";
        wait for Clk_period; 
        Features_din <= "0000000111010111";
        wait for Clk_period; 
        Features_din <= "1111101010001111";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000011111101";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110110111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001000010011";
        wait for Clk_period; 
        Features_din <= "0000000111110111";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000101011100";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "1111111001000000";
        wait for Clk_period; 
        Features_din <= "0000001000110101";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "0000001010100011";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "1111011100011010";
        wait for Clk_period; 
        Features_din <= "0000000011110011";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000001000111100";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000011000101";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001001100100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011100001";
        wait for Clk_period; 
        Features_din <= "0000001000111010";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "0000001011111100";
        wait for Clk_period; 
        Features_din <= "0000001001001110";
        wait for Clk_period; 
        Features_din <= "0000000110011110";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "1111111000110011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111011111001101";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110111110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "0000001001101100";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000001000101001";
        wait for Clk_period; 
        Features_din <= "0000000111110111";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000010100010111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "1111110100011001";
        wait for Clk_period; 
        Features_din <= "0000000101010111";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "1111100101100100";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "0000001000011011";
        wait for Clk_period; 
        Features_din <= "0000001100010010";
        wait for Clk_period; 
        Features_din <= "0000010100010001";
        wait for Clk_period; 
        Features_din <= "0000000101011001";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000001010001101";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000011011110";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001000001110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100000101";
        wait for Clk_period; 
        Features_din <= "0000001001001000";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000001100101001";
        wait for Clk_period; 
        Features_din <= "0000000111101110";
        wait for Clk_period; 
        Features_din <= "0000000111110110";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000010100011111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000100100010";
        wait for Clk_period; 
        Features_din <= "1111100011100010";
        wait for Clk_period; 
        Features_din <= "1111111000001110";
        wait for Clk_period; 
        Features_din <= "1111111010000011";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000000111100110";
        wait for Clk_period; 
        Features_din <= "0000001001000101";
        wait for Clk_period; 
        Features_din <= "0000010011011111";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111010101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "0000001000101101";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001000011100";
        wait for Clk_period; 
        Features_din <= "0000000111111001";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000000011010000";
        wait for Clk_period; 
        Features_din <= "1111101111111100";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000000011111101";
        wait for Clk_period; 
        Features_din <= "1111011111011100";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001010010101";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000001011110010";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000011100011";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001000000011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "1111111111101111";
        wait for Clk_period; 
        Features_din <= "0000001100000101";
        wait for Clk_period; 
        Features_din <= "0000000111010000";
        wait for Clk_period; 
        Features_din <= "0000000111000011";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000010001110100";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111110101110101";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111100010001011";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111010010000";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000001011011000";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010001110100";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000100110110";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001000001010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "0000001001010101";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "0000001100101100";
        wait for Clk_period; 
        Features_din <= "0000001000001101";
        wait for Clk_period; 
        Features_din <= "0000000111010010";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "1111110110110100";
        wait for Clk_period; 
        Features_din <= "0000000100001110";
        wait for Clk_period; 
        Features_din <= "0000000011101110";
        wait for Clk_period; 
        Features_din <= "0000000100000010";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "1111011110101111";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111110000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "0000001010001000";
        wait for Clk_period; 
        Features_din <= "1111111111100100";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000001000010110";
        wait for Clk_period; 
        Features_din <= "0000000111100101";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "1111100101000000";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000111000010";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "0000001010110000";
        wait for Clk_period; 
        Features_din <= "0000001000010111";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "1111101100100011";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000010101001100";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111001011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "0000001001111100";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "0000001100001110";
        wait for Clk_period; 
        Features_din <= "0000000111101011";
        wait for Clk_period; 
        Features_din <= "0000000110111011";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111100110101000";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000000110101010";
        wait for Clk_period; 
        Features_din <= "0000000100100111";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "0000000111100011";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000000101111001";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "1111101011101010";
        wait for Clk_period; 
        Features_din <= "0000001010110100";
        wait for Clk_period; 
        Features_din <= "0000010111010111";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000001011110011";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000101111111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011000011";
        wait for Clk_period; 
        Features_din <= "0000001001100100";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001000011000";
        wait for Clk_period; 
        Features_din <= "0000000111111100";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000001001101000";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "1111110001001011";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111011110101101";
        wait for Clk_period; 
        Features_din <= "0000001001101000";
        wait for Clk_period; 
        Features_din <= "0000001001101000";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000001001101000";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001001101000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000011100010";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111010001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "0000001000111100";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "0000001011111111";
        wait for Clk_period; 
        Features_din <= "0000000111111110";
        wait for Clk_period; 
        Features_din <= "0000000110111111";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111110101110100";
        wait for Clk_period; 
        Features_din <= "0000000101001001";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000001011111010";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "1111011111100010";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000010001100100";
        wait for Clk_period; 
        Features_din <= "0000001010011011";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000011000110";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001000101101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "0000001001010111";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000000111110101";
        wait for Clk_period; 
        Features_din <= "0000000111110101";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000010010111000";
        wait for Clk_period; 
        Features_din <= "0000001011110110";
        wait for Clk_period; 
        Features_din <= "1111110111100110";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "1111100011101011";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111000001111";
        wait for Clk_period; 
        Features_din <= "0000001001010111";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000011001001";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "0000010110001101";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000001010110001";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000011001100";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110101100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "0000001001001100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001000000000";
        wait for Clk_period; 
        Features_din <= "0000000111100100";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "1111100001011110";
        wait for Clk_period; 
        Features_din <= "1111110111100000";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "0000001001010110";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000011010000";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111001001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "0000001001111001";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000001000001111";
        wait for Clk_period; 
        Features_din <= "0000000111101000";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111101001111111";
        wait for Clk_period; 
        Features_din <= "0000001100110011";
        wait for Clk_period; 
        Features_din <= "0000010001111100";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000000111010010";
        wait for Clk_period; 
        Features_din <= "0000001000110100";
        wait for Clk_period; 
        Features_din <= "0000010011001010";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "1111110001101101";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111101111001010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000001001100011";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111011010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "0000001001010100";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "0000001100100010";
        wait for Clk_period; 
        Features_din <= "0000001000001010";
        wait for Clk_period; 
        Features_din <= "0000001000000010";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111110000001101";
        wait for Clk_period; 
        Features_din <= "0000000100101001";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001010110000";
        wait for Clk_period; 
        Features_din <= "0000000101011100";
        wait for Clk_period; 
        Features_din <= "0000000110010111";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000000011101111";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "1111110000111010";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "1111101001001001";
        wait for Clk_period; 
        Features_din <= "0000001001110110";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000110111010";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000011001001";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111011010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "0000001001001001";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000001100011010";
        wait for Clk_period; 
        Features_din <= "0000001001000110";
        wait for Clk_period; 
        Features_din <= "0000001000001101";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111101000101110";
        wait for Clk_period; 
        Features_din <= "0000001001010000";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000110111100";
        wait for Clk_period; 
        Features_din <= "0000001001100000";
        wait for Clk_period; 
        Features_din <= "0000001000011101";
        wait for Clk_period; 
        Features_din <= "1111111010000010";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "1111101101001111";
        wait for Clk_period; 
        Features_din <= "0000001010100101";
        wait for Clk_period; 
        Features_din <= "0000010111100101";
        wait for Clk_period; 
        Features_din <= "0000000100010000";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000111101010";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001010000110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011000100";
        wait for Clk_period; 
        Features_din <= "0000001000101111";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000001011110110";
        wait for Clk_period; 
        Features_din <= "0000001001001110";
        wait for Clk_period; 
        Features_din <= "0000000111001000";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "1111100100000010";
        wait for Clk_period; 
        Features_din <= "0000000011100000";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "1111101001100110";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000011100001";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001000000110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "0000001000110010";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "0000001100000101";
        wait for Clk_period; 
        Features_din <= "0000001001000100";
        wait for Clk_period; 
        Features_din <= "0000000111101011";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000010101110100";
        wait for Clk_period; 
        Features_din <= "0000000111100100";
        wait for Clk_period; 
        Features_din <= "0000000101010110";
        wait for Clk_period; 
        Features_din <= "0000000100110001";
        wait for Clk_period; 
        Features_din <= "0000000110010000";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "0000001010110100";
        wait for Clk_period; 
        Features_din <= "0000001000111001";
        wait for Clk_period; 
        Features_din <= "0000001000001010";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "1111101101100010";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "1111100100100111";
        wait for Clk_period; 
        Features_din <= "0000001011010011";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000101010110";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000011010111";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001000101100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "0000001001100000";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000001000010001";
        wait for Clk_period; 
        Features_din <= "0000000111010011";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000010100101001";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000001000111101";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000001001010101";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "0000001001011000";
        wait for Clk_period; 
        Features_din <= "0000001000110010";
        wait for Clk_period; 
        Features_din <= "0000001100100010";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "1111101011101001";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "1111100101011100";
        wait for Clk_period; 
        Features_din <= "0000000011011100";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111010100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "0000001000011111";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "0000001100110001";
        wait for Clk_period; 
        Features_din <= "0000001000110110";
        wait for Clk_period; 
        Features_din <= "0000000111111110";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "1111101010010111";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000000111011110";
        wait for Clk_period; 
        Features_din <= "0000001001000000";
        wait for Clk_period; 
        Features_din <= "0000000110000010";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001010111011";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "1111110011001110";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "1111101100110100";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000011010001";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111010111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "0000001001010101";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "0000001100011011";
        wait for Clk_period; 
        Features_din <= "0000001000010000";
        wait for Clk_period; 
        Features_din <= "0000000111101110";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000010100010001";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000001001110100";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "0000001100001000";
        wait for Clk_period; 
        Features_din <= "0000000111101000";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "1111101101111011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "1111100100111101";
        wait for Clk_period; 
        Features_din <= "0000001000001001";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000110111100";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000011011001";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110100101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000001100101100";
        wait for Clk_period; 
        Features_din <= "0000001000100010";
        wait for Clk_period; 
        Features_din <= "0000000111100000";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111100110001100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000001010100011";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "0000001001001101";
        wait for Clk_period; 
        Features_din <= "0000001000000001";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111101010110101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010100011000";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111010111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "0000001000101101";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "0000001100011110";
        wait for Clk_period; 
        Features_din <= "0000001001110010";
        wait for Clk_period; 
        Features_din <= "0000001000000001";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "1111101001111001";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000110011001";
        wait for Clk_period; 
        Features_din <= "0000000111010011";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111110011100001";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111101100110101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000000101000001";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111000101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "0000001001011010";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000001100001111";
        wait for Clk_period; 
        Features_din <= "0000001000111010";
        wait for Clk_period; 
        Features_din <= "0000000111011101";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000011011110010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111000101111";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "0000000011111101";
        wait for Clk_period; 
        Features_din <= "1111101111001111";
        wait for Clk_period; 
        Features_din <= "1111111001100111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111101101100111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111101001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "0000001100001110";
        wait for Clk_period; 
        Features_din <= "0000001001001101";
        wait for Clk_period; 
        Features_din <= "0000000110110100";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000000011001010";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "1111110110100100";
        wait for Clk_period; 
        Features_din <= "0000000100011011";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000011011011";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "1111011110110001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010001100000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010111101";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000011010110";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001000101111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100010010";
        wait for Clk_period; 
        Features_din <= "0000001000111100";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000001011110001";
        wait for Clk_period; 
        Features_din <= "0000001000000110";
        wait for Clk_period; 
        Features_din <= "0000000111000010";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111101000101110";
        wait for Clk_period; 
        Features_din <= "0000000101000100";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000000101001100";
        wait for Clk_period; 
        Features_din <= "0000010101101101";
        wait for Clk_period; 
        Features_din <= "0000000110101001";
        wait for Clk_period; 
        Features_din <= "0000000011011101";
        wait for Clk_period; 
        Features_din <= "0000000110010101";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "1111101010011110";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000001100000001";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000011000110";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001001111101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "0000001000101111";
        wait for Clk_period; 
        Features_din <= "1111111111111001";
        wait for Clk_period; 
        Features_din <= "0000001011101110";
        wait for Clk_period; 
        Features_din <= "0000001010101001";
        wait for Clk_period; 
        Features_din <= "0000000111010110";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000010101010010";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000000111111001";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "0000001011111001";
        wait for Clk_period; 
        Features_din <= "0000000101111011";
        wait for Clk_period; 
        Features_din <= "0000001011101100";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "1111101100000011";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "1111100110001011";
        wait for Clk_period; 
        Features_din <= "0000000111010011";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000100100010";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000011011101";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110111100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011100111";
        wait for Clk_period; 
        Features_din <= "0000001001111111";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000001100010110";
        wait for Clk_period; 
        Features_din <= "0000001001000111";
        wait for Clk_period; 
        Features_din <= "0000001000000001";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000010111011001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000110001100";
        wait for Clk_period; 
        Features_din <= "0000001001000000";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "0000000111111111";
        wait for Clk_period; 
        Features_din <= "0000001000110110";
        wait for Clk_period; 
        Features_din <= "0000000011001010";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "1111101100100111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "1111100101110010";
        wait for Clk_period; 
        Features_din <= "0000001100100110";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000111001010";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000011011100";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(2, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111000001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "0000001000100010";
        wait for Clk_period; 
        Features_din <= "1111111111100110";
        wait for Clk_period; 
        Features_din <= "0000001100100000";
        wait for Clk_period; 
        Features_din <= "0000000111111110";
        wait for Clk_period; 
        Features_din <= "0000001000010100";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111101010010011";
        wait for Clk_period; 
        Features_din <= "0000000110011100";
        wait for Clk_period; 
        Features_din <= "0000001100011100";
        wait for Clk_period; 
        Features_din <= "0000000100101010";
        wait for Clk_period; 
        Features_din <= "0000001011100000";
        wait for Clk_period; 
        Features_din <= "0000000110100011";
        wait for Clk_period; 
        Features_din <= "0000010001100011";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "1111110100001101";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "1111101100001010";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000010101101";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000100000111";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(3, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110111001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011001010";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000001100010010";
        wait for Clk_period; 
        Features_din <= "0000001000001001";
        wait for Clk_period; 
        Features_din <= "0000000111011010";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000010101011110";
        wait for Clk_period; 
        Features_din <= "0000000011010000";
        wait for Clk_period; 
        Features_din <= "0000001000100101";
        wait for Clk_period; 
        Features_din <= "0000000110110010";
        wait for Clk_period; 
        Features_din <= "0000001000000100";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "0000001001111001";
        wait for Clk_period; 
        Features_din <= "0000001000000100";
        wait for Clk_period; 
        Features_din <= "0000001100000011";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "1111101001001101";
        wait for Clk_period; 
        Features_din <= "0000000011110111";
        wait for Clk_period; 
        Features_din <= "1111101000000011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000100011001";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001000011011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011001000";
        wait for Clk_period; 
        Features_din <= "0000001000101100";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000001100010010";
        wait for Clk_period; 
        Features_din <= "0000001001001000";
        wait for Clk_period; 
        Features_din <= "0000000111000101";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "1111101000101000";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000101101100";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "0000001001110011";
        wait for Clk_period; 
        Features_din <= "0000001000001001";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111100111011011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000101000110";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110111001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "0000001001100011";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "0000001100010101";
        wait for Clk_period; 
        Features_din <= "0000000111011000";
        wait for Clk_period; 
        Features_din <= "0000000111010011";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111110101101110";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "1111100001010001";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000000110111011";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111110001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "0000001000110001";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000001100100111";
        wait for Clk_period; 
        Features_din <= "0000001000100001";
        wait for Clk_period; 
        Features_din <= "0000000111100000";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111101101000011";
        wait for Clk_period; 
        Features_din <= "0000000100011110";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000001001111011";
        wait for Clk_period; 
        Features_din <= "0000000101111110";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000000011111011";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "1111110001100100";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "1111101011100000";
        wait for Clk_period; 
        Features_din <= "0000001011111011";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000011101110";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(3, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110010000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011101101";
        wait for Clk_period; 
        Features_din <= "0000001001000111";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000001000100001";
        wait for Clk_period; 
        Features_din <= "0000001000011000";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000010100101101";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "1111110010000110";
        wait for Clk_period; 
        Features_din <= "0000000101010100";
        wait for Clk_period; 
        Features_din <= "0000001010101010";
        wait for Clk_period; 
        Features_din <= "1111101000100100";
        wait for Clk_period; 
        Features_din <= "1111110101101100";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "0000000111111100";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001010100101";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000000111001010";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000111010000";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000011100110";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001000010010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "0000001000110101";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000001100001010";
        wait for Clk_period; 
        Features_din <= "0000001000111000";
        wait for Clk_period; 
        Features_din <= "0000000111001011";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000010100111011";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000000111101011";
        wait for Clk_period; 
        Features_din <= "0000000110011110";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000001000011010";
        wait for Clk_period; 
        Features_din <= "0000001001110000";
        wait for Clk_period; 
        Features_din <= "0000000011111111";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "1111101100011011";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "1111100100101100";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000011011111";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111100010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011100110";
        wait for Clk_period; 
        Features_din <= "0000001001111011";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "0000001011110001";
        wait for Clk_period; 
        Features_din <= "0000001000101110";
        wait for Clk_period; 
        Features_din <= "0000000111001000";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000010100110000";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000001000000001";
        wait for Clk_period; 
        Features_din <= "0000000110000000";
        wait for Clk_period; 
        Features_din <= "0000000011110111";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "0000001010100111";
        wait for Clk_period; 
        Features_din <= "0000001000010000";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "1111101100100000";
        wait for Clk_period; 
        Features_din <= "0000001010001111";
        wait for Clk_period; 
        Features_din <= "1111100100111001";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000001100001110";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "0000000011101001";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111000010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "0000001001001010";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000001100001000";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000000111101110";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000000011101100";
        wait for Clk_period; 
        Features_din <= "0000000010111111";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111110101111111";
        wait for Clk_period; 
        Features_din <= "0000000101110011";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000001011000110";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "1111011110111110";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000001011000110";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000100010000";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111011000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011010010";
        wait for Clk_period; 
        Features_din <= "0000001001111111";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "0000001100000011";
        wait for Clk_period; 
        Features_din <= "0000001000011110";
        wait for Clk_period; 
        Features_din <= "0000000111011111";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000010011000000";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001011011000";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000000100100010";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "1111101011101001";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "1111100110111001";
        wait for Clk_period; 
        Features_din <= "0000000100010001";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000110111111";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000000011010011";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111001111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "0000001001001010";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000001100110001";
        wait for Clk_period; 
        Features_din <= "0000001000101111";
        wait for Clk_period; 
        Features_din <= "0000000111101101";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000010011001011";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "1111110010010111";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "1111100111000011";
        wait for Clk_period; 
        Features_din <= "1111110100110010";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "0000000101000101";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000001011000100";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000010011001011";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000011010110";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111000011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "0000001001011010";
        wait for Clk_period; 
        Features_din <= "1111111111101110";
        wait for Clk_period; 
        Features_din <= "0000001100000000";
        wait for Clk_period; 
        Features_din <= "0000001000111011";
        wait for Clk_period; 
        Features_din <= "0000000111001011";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111011100101100";
        wait for Clk_period; 
        Features_din <= "0000000101000011";
        wait for Clk_period; 
        Features_din <= "0000000100101111";
        wait for Clk_period; 
        Features_din <= "0000000011100010";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "1111111000110001";
        wait for Clk_period; 
        Features_din <= "0000000110011000";
        wait for Clk_period; 
        Features_din <= "0000000011000101";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000001011001001";
        wait for Clk_period; 
        Features_din <= "0000001011010010";
        wait for Clk_period; 
        Features_din <= "0000010001001101";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000001010001011";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000011010010";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110010011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "1111111111111010";
        wait for Clk_period; 
        Features_din <= "0000001100101011";
        wait for Clk_period; 
        Features_din <= "0000001000010101";
        wait for Clk_period; 
        Features_din <= "0000000111011100";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "1111110110100010";
        wait for Clk_period; 
        Features_din <= "0000000100110001";
        wait for Clk_period; 
        Features_din <= "0000000011101011";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "1111011110010101";
        wait for Clk_period; 
        Features_din <= "0000001001001000";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001000100110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "0000001011111010";
        wait for Clk_period; 
        Features_din <= "0000001000011100";
        wait for Clk_period; 
        Features_din <= "0000000111101110";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111011100000100";
        wait for Clk_period; 
        Features_din <= "0000001010101101";
        wait for Clk_period; 
        Features_din <= "0000001010110110";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "1111111001010101";
        wait for Clk_period; 
        Features_din <= "0000000110011110";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000010111101";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000001010111001";
        wait for Clk_period; 
        Features_din <= "0000001011011011";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001000001110";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000011001000";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110010101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100100000";
        wait for Clk_period; 
        Features_din <= "0000001001100011";
        wait for Clk_period; 
        Features_din <= "1111111111111011";
        wait for Clk_period; 
        Features_din <= "0000001100100011";
        wait for Clk_period; 
        Features_din <= "0000001000101100";
        wait for Clk_period; 
        Features_din <= "0000000111100111";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000010100111001";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "1111111001011000";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "1111100011100111";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111000100001";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "0000000101101110";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000010100000000";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000011100101";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111010101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "0000001001011100";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000001000010110";
        wait for Clk_period; 
        Features_din <= "0000000111110010";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111101100010101";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001000110111";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000101010101";
        wait for Clk_period; 
        Features_din <= "0000010010111011";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000000111001011";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "1111110011000100";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "1111101011010011";
        wait for Clk_period; 
        Features_din <= "0000001011001010";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000011101110";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000011101110";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001000011111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "0000001000010000";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "0000001001010100";
        wait for Clk_period; 
        Features_din <= "0000000110110100";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "1111101010000011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001011011001";
        wait for Clk_period; 
        Features_din <= "0000001010110001";
        wait for Clk_period; 
        Features_din <= "0000000110010001";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010010100001";
        wait for Clk_period; 
        Features_din <= "0000000011001100";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "1111110100010011";
        wait for Clk_period; 
        Features_din <= "0000000011011110";
        wait for Clk_period; 
        Features_din <= "1111101100011011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000011010101";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111110011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011001111";
        wait for Clk_period; 
        Features_din <= "0000001001111000";
        wait for Clk_period; 
        Features_din <= "1111111111110110";
        wait for Clk_period; 
        Features_din <= "0000001100010001";
        wait for Clk_period; 
        Features_din <= "0000001001111111";
        wait for Clk_period; 
        Features_din <= "0000000111011001";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111101010011011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000000111100101";
        wait for Clk_period; 
        Features_din <= "0000000101001010";
        wait for Clk_period; 
        Features_din <= "0000000101011101";
        wait for Clk_period; 
        Features_din <= "0000010010000100";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "1111110011001110";
        wait for Clk_period; 
        Features_din <= "0000000111111010";
        wait for Clk_period; 
        Features_din <= "1111101101000001";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110101010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000001000100010";
        wait for Clk_period; 
        Features_din <= "0000000111111101";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "1111101010111011";
        wait for Clk_period; 
        Features_din <= "0000000111101001";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000000100101000";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000000110100111";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000001011100101";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "1111110011001011";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "1111101100001011";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111101100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "0000001000111101";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000001100100011";
        wait for Clk_period; 
        Features_din <= "0000001000011101";
        wait for Clk_period; 
        Features_din <= "0000000111111010";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "1111100101011011";
        wait for Clk_period; 
        Features_din <= "0000000101110011";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "1111101000000010";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000011001101";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111110011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011011010";
        wait for Clk_period; 
        Features_din <= "0000001010000001";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "0000001100001111";
        wait for Clk_period; 
        Features_din <= "0000001000001111";
        wait for Clk_period; 
        Features_din <= "0000000111010010";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111011011001110";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000000111100111";
        wait for Clk_period; 
        Features_din <= "0000000111111111";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "0000001000000010";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000011000010";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "0000001010011110";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000111111110";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000011010111";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110011000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "0000001001010011";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000001100010111";
        wait for Clk_period; 
        Features_din <= "0000001001000110";
        wait for Clk_period; 
        Features_din <= "0000000111111101";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000000110011000";
        wait for Clk_period; 
        Features_din <= "0000000011101111";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "1111110110011100";
        wait for Clk_period; 
        Features_din <= "0000000100011100";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000001011110010";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "1111011110001111";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000100101111";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111000010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011101110";
        wait for Clk_period; 
        Features_din <= "0000001001011100";
        wait for Clk_period; 
        Features_din <= "1111111111111110";
        wait for Clk_period; 
        Features_din <= "0000001100100100";
        wait for Clk_period; 
        Features_din <= "0000001000001111";
        wait for Clk_period; 
        Features_din <= "0000000111101111";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111101100101000";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "0000000111110001";
        wait for Clk_period; 
        Features_din <= "0000001001111111";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "1111110010101110";
        wait for Clk_period; 
        Features_din <= "1111110110000001";
        wait for Clk_period; 
        Features_din <= "0000001001110011";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000010001110001";
        wait for Clk_period; 
        Features_din <= "0000000101000010";
        wait for Clk_period; 
        Features_din <= "0000011100011100";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000001011101011";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000011011011";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001000110010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011000010";
        wait for Clk_period; 
        Features_din <= "0000001001010101";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "0000001100101010";
        wait for Clk_period; 
        Features_din <= "0000001000101000";
        wait for Clk_period; 
        Features_din <= "0000000111111110";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111101011000100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000000110110110";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000101110101";
        wait for Clk_period; 
        Features_din <= "0000010001111111";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001010101110";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "1111110011100001";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "1111101011111111";
        wait for Clk_period; 
        Features_din <= "0000001001011011";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000011000010";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "0000000011110111";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110010100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "0000001001101000";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "0000001101000100";
        wait for Clk_period; 
        Features_din <= "0000001001000010";
        wait for Clk_period; 
        Features_din <= "0000001000000011";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111101111111000";
        wait for Clk_period; 
        Features_din <= "0000001100100011";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001000101011";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "0000000011011110";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "0000011110000001";
        wait for Clk_period; 
        Features_din <= "0000000100010000";
        wait for Clk_period; 
        Features_din <= "1111101100100010";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000001000111111";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000011100010";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110110001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "0000001000110000";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000001100011011";
        wait for Clk_period; 
        Features_din <= "0000001000010011";
        wait for Clk_period; 
        Features_din <= "0000000111101001";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "1111011110010100";
        wait for Clk_period; 
        Features_din <= "0000000101000010";
        wait for Clk_period; 
        Features_din <= "0000000110101001";
        wait for Clk_period; 
        Features_din <= "0000001001000100";
        wait for Clk_period; 
        Features_din <= "0000000101011001";
        wait for Clk_period; 
        Features_din <= "1111110110110010";
        wait for Clk_period; 
        Features_din <= "0000001010010011";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "0000000010111111";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000001000000111";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010010110110";
        wait for Clk_period; 
        Features_din <= "0000001011101010";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000110100100";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000010111110";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111001110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011111001";
        wait for Clk_period; 
        Features_din <= "0000001000111010";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001000011011";
        wait for Clk_period; 
        Features_din <= "0000001000010110";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "1111101001001011";
        wait for Clk_period; 
        Features_din <= "0000000010101100";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "1111100100011001";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001001110010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010011100";
        wait for Clk_period; 
        Features_din <= "0000001001011011";
        wait for Clk_period; 
        Features_din <= "1111111111011011";
        wait for Clk_period; 
        Features_din <= "0000001011101111";
        wait for Clk_period; 
        Features_din <= "0000001001010110";
        wait for Clk_period; 
        Features_din <= "0000000110101011";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001000111100";
        wait for Clk_period; 
        Features_din <= "0000000011101101";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "1111110110001110";
        wait for Clk_period; 
        Features_din <= "1111100010010100";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "0000000110000011";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000010101101010";
        wait for Clk_period; 
        Features_din <= "0000000011000010";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000110110000";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001001001110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011111111";
        wait for Clk_period; 
        Features_din <= "0000001000100101";
        wait for Clk_period; 
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "0000001000111000";
        wait for Clk_period; 
        Features_din <= "0000000111000110";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111101100101111";
        wait for Clk_period; 
        Features_din <= "0000000110100111";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000000101000110";
        wait for Clk_period; 
        Features_din <= "0000000110000001";
        wait for Clk_period; 
        Features_din <= "0000000111010000";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "1111110010110100";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "1111101010011100";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000110110000";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001000010111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000001100010010";
        wait for Clk_period; 
        Features_din <= "0000001000101111";
        wait for Clk_period; 
        Features_din <= "0000000111101001";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "1111101000110001";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000001010011011";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000011101111";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000001001010010";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "1111100110100001";
        wait for Clk_period; 
        Features_din <= "0000000100100011";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000011010000";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110110100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "0000001001100011";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000001100011110";
        wait for Clk_period; 
        Features_din <= "0000001001001010";
        wait for Clk_period; 
        Features_din <= "0000000111110111";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000010111011100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000110111100";
        wait for Clk_period; 
        Features_din <= "0000000011111100";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "0000001001001101";
        wait for Clk_period; 
        Features_din <= "0000000111101011";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "1111101100100110";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "1111100110000111";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000011111011";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000011011110";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110011001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "0000001001111100";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000001000000111";
        wait for Clk_period; 
        Features_din <= "0000001000000101";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000010100010101";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000100001010";
        wait for Clk_period; 
        Features_din <= "0000001001000100";
        wait for Clk_period; 
        Features_din <= "1111111001101000";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "0000000110010100";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000001010111010";
        wait for Clk_period; 
        Features_din <= "0000000101011001";
        wait for Clk_period; 
        Features_din <= "1111011101101111";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110001100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "0000001001011100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000001000111100";
        wait for Clk_period; 
        Features_din <= "0000001000000000";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000001100111000";
        wait for Clk_period; 
        Features_din <= "0000001000100011";
        wait for Clk_period; 
        Features_din <= "1111111010101010";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000001001011101";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111100100001010";
        wait for Clk_period; 
        Features_din <= "0000001100100000";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "0000010101001010";
        wait for Clk_period; 
        Features_din <= "0000000100001000";
        wait for Clk_period; 
        Features_din <= "1111110001010010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000000010111100";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000001100111000";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000100010000";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110001111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011101010";
        wait for Clk_period; 
        Features_din <= "0000001001000011";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001000100101";
        wait for Clk_period; 
        Features_din <= "0000000111010100";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000010011001011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111000111100";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111100010010100";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111010000100";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000001000100010";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010011001011";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000100001111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111001110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "0000001001101000";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "0000001100010110";
        wait for Clk_period; 
        Features_din <= "0000001001000100";
        wait for Clk_period; 
        Features_din <= "0000000111110110";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000010001110010";
        wait for Clk_period; 
        Features_din <= "0000000101001100";
        wait for Clk_period; 
        Features_din <= "0000001011001010";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "0000001011101100";
        wait for Clk_period; 
        Features_din <= "0000000110111101";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "1111101101101110";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111100011001010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110101111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "0000001010010101";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "0000001100001000";
        wait for Clk_period; 
        Features_din <= "0000001000111110";
        wait for Clk_period; 
        Features_din <= "0000000111111110";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000010100111001";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000001000111101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "0000001010011001";
        wait for Clk_period; 
        Features_din <= "0000000111101101";
        wait for Clk_period; 
        Features_din <= "0000000111010100";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "1111101011101111";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "1111100101100111";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001010010001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010100110";
        wait for Clk_period; 
        Features_din <= "0000001000110011";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "0000001100001010";
        wait for Clk_period; 
        Features_din <= "0000000111111001";
        wait for Clk_period; 
        Features_din <= "0000000111001011";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111101111101010";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000011101101110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101100011110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000011001101";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111011110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "0000001001101010";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "0000001100000000";
        wait for Clk_period; 
        Features_din <= "0000001001101001";
        wait for Clk_period; 
        Features_din <= "0000000111011010";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000010001111100";
        wait for Clk_period; 
        Features_din <= "0000000100101101";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "0000000011100110";
        wait for Clk_period; 
        Features_din <= "0000000100011001";
        wait for Clk_period; 
        Features_din <= "1111110100111010";
        wait for Clk_period; 
        Features_din <= "0000001000101111";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "1111011111110111";
        wait for Clk_period; 
        Features_din <= "0000001010111110";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000001010101010";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000011010000";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111110010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011111101";
        wait for Clk_period; 
        Features_din <= "0000001001000011";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000001001011010";
        wait for Clk_period; 
        Features_din <= "0000001000000010";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000010010101000";
        wait for Clk_period; 
        Features_din <= "0000000101110000";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000000100001000";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "0000000110100011";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "1111101010111110";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "1111100111100011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111001111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100010111";
        wait for Clk_period; 
        Features_din <= "0000001001010100";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000001100101001";
        wait for Clk_period; 
        Features_din <= "0000001000101111";
        wait for Clk_period; 
        Features_din <= "0000000111101111";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "1111110110001000";
        wait for Clk_period; 
        Features_din <= "0000000101100000";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "1111011110110001";
        wait for Clk_period; 
        Features_din <= "0000001010011011";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000001100000110";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111011001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "0000001001001000";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "0000001100001110";
        wait for Clk_period; 
        Features_din <= "0000001000101011";
        wait for Clk_period; 
        Features_din <= "0000001000010100";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000011001000011";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "1111111001001000";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000001000011111";
        wait for Clk_period; 
        Features_din <= "1111100100111111";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111000010111";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "0000000100101101";
        wait for Clk_period; 
        Features_din <= "0000000110011110";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110011000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000001100011011";
        wait for Clk_period; 
        Features_din <= "0000001000000110";
        wait for Clk_period; 
        Features_din <= "0000000111101111";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000010010100000";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "0000000111011010";
        wait for Clk_period; 
        Features_din <= "0000001001001011";
        wait for Clk_period; 
        Features_din <= "0000001000011000";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000000110011100";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "1111110001000001";
        wait for Clk_period; 
        Features_din <= "0000001000110101";
        wait for Clk_period; 
        Features_din <= "1111100001011010";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000001101000100";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000010111101";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111100110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "0000001001111100";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000001100011001";
        wait for Clk_period; 
        Features_din <= "0000001000101100";
        wait for Clk_period; 
        Features_din <= "0000000111011011";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111100111111010";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000001000101101";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000001100010011";
        wait for Clk_period; 
        Features_din <= "0000001010011010";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "1111100111001100";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000011001010";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110111110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100000001";
        wait for Clk_period; 
        Features_din <= "0000001001101101";
        wait for Clk_period; 
        Features_din <= "1111111111111000";
        wait for Clk_period; 
        Features_din <= "0000001100010000";
        wait for Clk_period; 
        Features_din <= "0000001001000100";
        wait for Clk_period; 
        Features_din <= "0000000111111001";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "1111101110001101";
        wait for Clk_period; 
        Features_din <= "0000000011100110";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001011001000";
        wait for Clk_period; 
        Features_din <= "0000000100111101";
        wait for Clk_period; 
        Features_din <= "0000000011101000";
        wait for Clk_period; 
        Features_din <= "0000010011111101";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000001001111011";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "1111110101000011";
        wait for Clk_period; 
        Features_din <= "0000001011110101";
        wait for Clk_period; 
        Features_din <= "1111101000110010";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000001010001010";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000011101001";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111110010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "0000001001000101";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000001100101010";
        wait for Clk_period; 
        Features_din <= "0000001001000000";
        wait for Clk_period; 
        Features_din <= "0000000111011110";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "1111100110100111";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "0000001001101010";
        wait for Clk_period; 
        Features_din <= "0000000110010111";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "1111101010110110";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000110110111";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000011000111";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001001001010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011010101";
        wait for Clk_period; 
        Features_din <= "0000001001011010";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000001100010111";
        wait for Clk_period; 
        Features_din <= "0000001000101000";
        wait for Clk_period; 
        Features_din <= "0000000111011011";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000010100000010";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "1111110101111111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "1111100100011011";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111000100101";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000001011011010";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000010010000001";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000010111101";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110111010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100001100";
        wait for Clk_period; 
        Features_din <= "0000001001000111";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001000100010";
        wait for Clk_period; 
        Features_din <= "0000000111010011";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "1111101100110001";
        wait for Clk_period; 
        Features_din <= "0000000110100110";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "0000001010101100";
        wait for Clk_period; 
        Features_din <= "0000000101110100";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001011011100";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "1111110010000000";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111101011011010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110110110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "0000001001100011";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000001100011000";
        wait for Clk_period; 
        Features_din <= "0000001000011011";
        wait for Clk_period; 
        Features_din <= "0000000111001100";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000010001101101";
        wait for Clk_period; 
        Features_din <= "0000000111001101";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "1111100001011100";
        wait for Clk_period; 
        Features_din <= "1111111001011010";
        wait for Clk_period; 
        Features_din <= "1111110110010101";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000001001010110";
        wait for Clk_period; 
        Features_din <= "0000001000000111";
        wait for Clk_period; 
        Features_din <= "0000010001110001";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000001011110001";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000010110011";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001000111001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000001011111111";
        wait for Clk_period; 
        Features_din <= "0000001000100111";
        wait for Clk_period; 
        Features_din <= "0000000111110011";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000010011000100";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001011001110";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "0000001010010000";
        wait for Clk_period; 
        Features_din <= "0000000111110110";
        wait for Clk_period; 
        Features_din <= "0000000111100111";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "1111101001011111";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111100110111011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000110100100";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000011100100";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110011101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100001001";
        wait for Clk_period; 
        Features_din <= "0000001001010101";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000001000010010";
        wait for Clk_period; 
        Features_din <= "0000000111100110";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "1111011110111000";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000001011101011";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000000110001101";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000111110000";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110000001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100001000";
        wait for Clk_period; 
        Features_din <= "0000001000101111";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000000111110100";
        wait for Clk_period; 
        Features_din <= "0000001000001000";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111011011001010";
        wait for Clk_period; 
        Features_din <= "0000000101000011";
        wait for Clk_period; 
        Features_din <= "0000000111011001";
        wait for Clk_period; 
        Features_din <= "0000001100101000";
        wait for Clk_period; 
        Features_din <= "0000000111100100";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "0000000101001011";
        wait for Clk_period; 
        Features_din <= "0000000110010011";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000001011011000";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001001001011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "0000001001101100";
        wait for Clk_period; 
        Features_din <= "1111111111110101";
        wait for Clk_period; 
        Features_din <= "0000001100001011";
        wait for Clk_period; 
        Features_din <= "0000001000110111";
        wait for Clk_period; 
        Features_din <= "0000000110101011";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111100101100101";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "0000001011000110";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000000101101101";
        wait for Clk_period; 
        Features_din <= "0000001011001111";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "1111101011101101";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000010010110011";
        wait for Clk_period; 
        Features_din <= "0000001010111010";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000011111000";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000011010001";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111011111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "0000001001100011";
        wait for Clk_period; 
        Features_din <= "1111111111110010";
        wait for Clk_period; 
        Features_din <= "0000001100010001";
        wait for Clk_period; 
        Features_din <= "0000001000110000";
        wait for Clk_period; 
        Features_din <= "0000000111011110";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000010100001001";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "0000001000101000";
        wait for Clk_period; 
        Features_din <= "0000000010111100";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000000110010110";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "1111101100000100";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "1111100101011100";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000011001110";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001001000101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "0000001000011100";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "0000001100011101";
        wait for Clk_period; 
        Features_din <= "0000001001011011";
        wait for Clk_period; 
        Features_din <= "0000000111011100";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111101011111111";
        wait for Clk_period; 
        Features_din <= "0000001001110001";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000001001110100";
        wait for Clk_period; 
        Features_din <= "0000000101100101";
        wait for Clk_period; 
        Features_din <= "0000010011011001";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001100101001";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "1111110011101000";
        wait for Clk_period; 
        Features_din <= "0000001001001100";
        wait for Clk_period; 
        Features_din <= "1111101011001101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000001000101111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111101111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011010011";
        wait for Clk_period; 
        Features_din <= "0000001001000111";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        Features_din <= "0000001001010101";
        wait for Clk_period; 
        Features_din <= "0000000111100010";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000010011000111";
        wait for Clk_period; 
        Features_din <= "0000000110010000";
        wait for Clk_period; 
        Features_din <= "0000001010101100";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "0000001011101111";
        wait for Clk_period; 
        Features_din <= "0000000110101110";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "1111101100001001";
        wait for Clk_period; 
        Features_din <= "0000001010000000";
        wait for Clk_period; 
        Features_din <= "1111100100111011";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000001010110100";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111001011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "0000001001000101";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000001100100000";
        wait for Clk_period; 
        Features_din <= "0000001000110000";
        wait for Clk_period; 
        Features_din <= "0000000111011011";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001011010000";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000000100011001";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "1111101010001101";
        wait for Clk_period; 
        Features_din <= "0000000100111011";
        wait for Clk_period; 
        Features_din <= "1111100111001110";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000001010010000";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111001010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011101011";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001001000000";
        wait for Clk_period; 
        Features_din <= "0000000111101011";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111100111110101";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000000101001000";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "1111110111010010";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000011011001110";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "1111110010001100";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000101001100";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000011001110";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110000110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100100110";
        wait for Clk_period; 
        Features_din <= "0000001001011111";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000000111110111";
        wait for Clk_period; 
        Features_din <= "0000001000011101";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000010110000111";
        wait for Clk_period; 
        Features_din <= "0000001010000001";
        wait for Clk_period; 
        Features_din <= "1111111000101000";
        wait for Clk_period; 
        Features_din <= "0000000011101011";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "1111100011100110";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111001101010";
        wait for Clk_period; 
        Features_din <= "0000000101010000";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000100111001";
        wait for Clk_period; 
        Features_din <= "0000001001110100";
        wait for Clk_period; 
        Features_din <= "0000010011000010";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000111101110";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000011010010";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110110110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011100011";
        wait for Clk_period; 
        Features_din <= "0000001001110000";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "0000001100011010";
        wait for Clk_period; 
        Features_din <= "0000001001101000";
        wait for Clk_period; 
        Features_din <= "0000000111100110";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111011100101111";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000100100011";
        wait for Clk_period; 
        Features_din <= "0000000100100011";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "1111111000110100";
        wait for Clk_period; 
        Features_din <= "0000000110101000";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000001010001000";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111110010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "0000001000110011";
        wait for Clk_period; 
        Features_din <= "1111111111101010";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001000101110";
        wait for Clk_period; 
        Features_din <= "0000001000010000";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111100110000100";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000000011111000";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "1111110111001110";
        wait for Clk_period; 
        Features_din <= "0000001011110001";
        wait for Clk_period; 
        Features_din <= "1111101110100001";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000000111110100";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000010001110011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000100001110";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000011001010";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001000111101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000001100011000";
        wait for Clk_period; 
        Features_din <= "0000001000011000";
        wait for Clk_period; 
        Features_din <= "0000000111010011";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000000110010011";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000110110000";
        wait for Clk_period; 
        Features_din <= "1111110110010001";
        wait for Clk_period; 
        Features_din <= "0000000011101000";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "1111011111000101";
        wait for Clk_period; 
        Features_din <= "0000001011000011";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000011010001";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(3, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110011100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "0000001001000111";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000001100011100";
        wait for Clk_period; 
        Features_din <= "0000001000100010";
        wait for Clk_period; 
        Features_din <= "0000000111101011";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000110010000";
        wait for Clk_period; 
        Features_din <= "0000000100111000";
        wait for Clk_period; 
        Features_din <= "0000011110111010";
        wait for Clk_period; 
        Features_din <= "0000001100101100";
        wait for Clk_period; 
        Features_din <= "0000000100011000";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "0000000011010011";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "1111100100110011";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "0000001000000101";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000101110101";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000100100001";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(2, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110001000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "0000001001101000";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000000111101110";
        wait for Clk_period; 
        Features_din <= "0000000111111000";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111101100101010";
        wait for Clk_period; 
        Features_din <= "0000000101100000";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000000110010010";
        wait for Clk_period; 
        Features_din <= "0000000110010110";
        wait for Clk_period; 
        Features_din <= "0000000101111110";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111110000001100";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "1111101101000101";
        wait for Clk_period; 
        Features_din <= "0000001000101001";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000111011100";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000011111110";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001011001010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010010000";
        wait for Clk_period; 
        Features_din <= "0000001000111000";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "0000001100000000";
        wait for Clk_period; 
        Features_din <= "0000001001010010";
        wait for Clk_period; 
        Features_din <= "0000000111001011";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000010110110110";
        wait for Clk_period; 
        Features_din <= "0000000101010101";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "0000001000000001";
        wait for Clk_period; 
        Features_din <= "0000001100010100";
        wait for Clk_period; 
        Features_din <= "0000000110101110";
        wait for Clk_period; 
        Features_din <= "1111110100111110";
        wait for Clk_period; 
        Features_din <= "1111110101111111";
        wait for Clk_period; 
        Features_din <= "0000000110010110";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000010100011010";
        wait for Clk_period; 
        Features_din <= "0000001100001101";
        wait for Clk_period; 
        Features_din <= "1111101000010111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000001000111000";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000010111111";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001010001101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011011001";
        wait for Clk_period; 
        Features_din <= "0000001000111000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000001011001111";
        wait for Clk_period; 
        Features_din <= "0000001000101000";
        wait for Clk_period; 
        Features_din <= "0000000110011011";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111110000111001";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000011101111110";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "1111101100000010";
        wait for Clk_period; 
        Features_din <= "0000000110101110";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000101101111";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000011010111";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001001000010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011010000";
        wait for Clk_period; 
        Features_din <= "0000001001010000";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "0000001000011110";
        wait for Clk_period; 
        Features_din <= "0000000111000110";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000010100111101";
        wait for Clk_period; 
        Features_din <= "0000000110000000";
        wait for Clk_period; 
        Features_din <= "0000000111010110";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000111001101";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "0000001011011010";
        wait for Clk_period; 
        Features_din <= "0000001000000000";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "1111101100101011";
        wait for Clk_period; 
        Features_din <= "0000000011000101";
        wait for Clk_period; 
        Features_din <= "1111100100111111";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000011001111";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001000000100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011010111";
        wait for Clk_period; 
        Features_din <= "0000001000011110";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000001000111100";
        wait for Clk_period; 
        Features_din <= "0000001000010100";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000001011000111";
        wait for Clk_period; 
        Features_din <= "0000000100000110";
        wait for Clk_period; 
        Features_din <= "0000001011010100";
        wait for Clk_period; 
        Features_din <= "0000000110010010";
        wait for Clk_period; 
        Features_din <= "0000000110001101";
        wait for Clk_period; 
        Features_din <= "1111110111110000";
        wait for Clk_period; 
        Features_din <= "0000000110011001";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "1111011101010111";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000000100000010";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000110101000";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000010111110";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111000001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011011000";
        wait for Clk_period; 
        Features_din <= "0000001001000111";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000001000111111";
        wait for Clk_period; 
        Features_din <= "0000000111011010";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111110110000000";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000100110000000";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "1111111000001000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "1111110110000101";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "1111111000001000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000111000000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "0000001001000101";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "0000001001001011";
        wait for Clk_period; 
        Features_din <= "0000001000011000";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111101000011100";
        wait for Clk_period; 
        Features_din <= "0000000111010101";
        wait for Clk_period; 
        Features_din <= "0000001010100011";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000001010100000";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000001100010000";
        wait for Clk_period; 
        Features_din <= "0000001000111011";
        wait for Clk_period; 
        Features_din <= "0000001100000100";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111100111000111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000010111000";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110110001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "0000001000010110";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000001001101001";
        wait for Clk_period; 
        Features_din <= "0000000111000010";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000011000010001";
        wait for Clk_period; 
        Features_din <= "0000000011011100";
        wait for Clk_period; 
        Features_din <= "0000000111001001";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000001100010000";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "0000001000111011";
        wait for Clk_period; 
        Features_din <= "0000000110100110";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "1111101100100101";
        wait for Clk_period; 
        Features_din <= "0000001011010010";
        wait for Clk_period; 
        Features_din <= "1111100110100011";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000001010110100";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
            wait;
    end process;
end;
